library work;
use work.keccak_globals.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rho_pi_chi is
    port(
        rho_pi_chi_in : in k_state;
        rho_pi_chi_out: out k_state
    );
end entity rho_pi_chi;

architecture RTL of rho_pi_chi is

    signal pi_in,pi_out,rho_in,rho_out,chi_in,chi_out : k_state;


begin

    rho_in <= rho_pi_chi_in;
    ----------------------------
    --rho_1-----------------------
    ----------------------------
    i4001: for i in 0 to 63 generate
        rho_out(0)(0)(i)<=rho_in(0)(0)(i);
    end generate;
    i4002: for i in 0 to 63 generate
        rho_out(0)(1)(i)<=rho_in(0)(1)((i-1)mod 64);
    end generate;
    i4003: for i in 0 to 63 generate
        rho_out(0)(2)(i)<=rho_in(0)(2)((i-62)mod 64);
    end generate;
    i4004: for i in 0 to 63 generate
        rho_out(0)(3)(i)<=rho_in(0)(3)((i-28)mod 64);
    end generate;
    i4005: for i in 0 to 63 generate
        rho_out(0)(4)(i)<=rho_in(0)(4)((i-27)mod 64);
    end generate;

    i4011: for i in 0 to 63 generate
        rho_out(1)(0)(i)<=rho_in(1)(0)((i-36)mod 64);
    end generate;
    i4012: for i in 0 to 63 generate
        rho_out(1)(1)(i)<=rho_in(1)(1)((i-44)mod 64);
    end generate;
    i4013: for i in 0 to 63 generate
        rho_out(1)(2)(i)<=rho_in(1)(2)((i-6)mod 64);
    end generate;
    i4014: for i in 0 to 63 generate
        rho_out(1)(3)(i)<=rho_in(1)(3)((i-55)mod 64);
    end generate;
    i4015: for i in 0 to 63 generate
        rho_out(1)(4)(i)<=rho_in(1)(4)((i-20)mod 64);
    end generate;

    i4021: for i in 0 to 63 generate
        rho_out(2)(0)(i)<=rho_in(2)(0)((i-3)mod 64);
    end generate;
    i4022: for i in 0 to 63 generate
        rho_out(2)(1)(i)<=rho_in(2)(1)((i-10)mod 64);
    end generate;
    i4023: for i in 0 to 63 generate
        rho_out(2)(2)(i)<=rho_in(2)(2)((i-43)mod 64);
    end generate;
    i4024: for i in 0 to 63 generate
        rho_out(2)(3)(i)<=rho_in(2)(3)((i-25)mod 64);
    end generate;
    i4025: for i in 0 to 63 generate
        rho_out(2)(4)(i)<=rho_in(2)(4)((i-39)mod 64);
    end generate;

    i4031: for i in 0 to 63 generate
        rho_out(3)(0)(i)<=rho_in(3)(0)((i-41)mod 64);
    end generate;
    i4032: for i in 0 to 63 generate
        rho_out(3)(1)(i)<=rho_in(3)(1)((i-45)mod 64);
    end generate;
    i4033: for i in 0 to 63 generate
        rho_out(3)(2)(i)<=rho_in(3)(2)((i-15)mod 64);
    end generate;
    i4034: for i in 0 to 63 generate
        rho_out(3)(3)(i)<=rho_in(3)(3)((i-21)mod 64);
    end generate;
    i4035: for i in 0 to 63 generate
        rho_out(3)(4)(i)<=rho_in(3)(4)((i-8)mod 64);
    end generate;

    i4041: for i in 0 to 63 generate
        rho_out(4)(0)(i)<=rho_in(4)(0)((i-18)mod 64);
    end generate;
    i4042: for i in 0 to 63 generate
        rho_out(4)(1)(i)<=rho_in(4)(1)((i-2)mod 64);
    end generate;
    i4043: for i in 0 to 63 generate
        rho_out(4)(2)(i)<=rho_in(4)(2)((i-61)mod 64);
    end generate;
    i4044: for i in 0 to 63 generate
        rho_out(4)(3)(i)<=rho_in(4)(3)((i-56)mod 64);
    end generate;
    i4045: for i in 0 to 63 generate
        rho_out(4)(4)(i)<=rho_in(4)(4)((i-14)mod 64);
    end generate;


    pi_in <= rho_out;
    -------------------------
    -- pi + chi  -----------------
    -------------------------



    

chi_out(0)(0)(0) <= pi_in(0)(0)(0) xor ((not pi_in(1)(1)(0)) and pi_in(2)(2)(0));
 chi_out(0)(0)(1) <= pi_in(0)(0)(1) xor ((not pi_in(1)(1)(1)) and pi_in(2)(2)(1));
 chi_out(0)(0)(2) <= pi_in(0)(0)(2) xor ((not pi_in(1)(1)(2)) and pi_in(2)(2)(2));
 chi_out(0)(0)(3) <= pi_in(0)(0)(3) xor ((not pi_in(1)(1)(3)) and pi_in(2)(2)(3));
 chi_out(0)(0)(4) <= pi_in(0)(0)(4) xor ((not pi_in(1)(1)(4)) and pi_in(2)(2)(4));
 chi_out(0)(0)(5) <= pi_in(0)(0)(5) xor ((not pi_in(1)(1)(5)) and pi_in(2)(2)(5));
 chi_out(0)(0)(6) <= pi_in(0)(0)(6) xor ((not pi_in(1)(1)(6)) and pi_in(2)(2)(6));
 chi_out(0)(0)(7) <= pi_in(0)(0)(7) xor ((not pi_in(1)(1)(7)) and pi_in(2)(2)(7));
 chi_out(0)(0)(8) <= pi_in(0)(0)(8) xor ((not pi_in(1)(1)(8)) and pi_in(2)(2)(8));
 chi_out(0)(0)(9) <= pi_in(0)(0)(9) xor ((not pi_in(1)(1)(9)) and pi_in(2)(2)(9));
 chi_out(0)(0)(10) <= pi_in(0)(0)(10) xor ((not pi_in(1)(1)(10)) and pi_in(2)(2)(10));
 chi_out(0)(0)(11) <= pi_in(0)(0)(11) xor ((not pi_in(1)(1)(11)) and pi_in(2)(2)(11));
 chi_out(0)(0)(12) <= pi_in(0)(0)(12) xor ((not pi_in(1)(1)(12)) and pi_in(2)(2)(12));
 chi_out(0)(0)(13) <= pi_in(0)(0)(13) xor ((not pi_in(1)(1)(13)) and pi_in(2)(2)(13));
 chi_out(0)(0)(14) <= pi_in(0)(0)(14) xor ((not pi_in(1)(1)(14)) and pi_in(2)(2)(14));
 chi_out(0)(0)(15) <= pi_in(0)(0)(15) xor ((not pi_in(1)(1)(15)) and pi_in(2)(2)(15));
 chi_out(0)(0)(16) <= pi_in(0)(0)(16) xor ((not pi_in(1)(1)(16)) and pi_in(2)(2)(16));
 chi_out(0)(0)(17) <= pi_in(0)(0)(17) xor ((not pi_in(1)(1)(17)) and pi_in(2)(2)(17));
 chi_out(0)(0)(18) <= pi_in(0)(0)(18) xor ((not pi_in(1)(1)(18)) and pi_in(2)(2)(18));
 chi_out(0)(0)(19) <= pi_in(0)(0)(19) xor ((not pi_in(1)(1)(19)) and pi_in(2)(2)(19));
 chi_out(0)(0)(20) <= pi_in(0)(0)(20) xor ((not pi_in(1)(1)(20)) and pi_in(2)(2)(20));
 chi_out(0)(0)(21) <= pi_in(0)(0)(21) xor ((not pi_in(1)(1)(21)) and pi_in(2)(2)(21));
 chi_out(0)(0)(22) <= pi_in(0)(0)(22) xor ((not pi_in(1)(1)(22)) and pi_in(2)(2)(22));
 chi_out(0)(0)(23) <= pi_in(0)(0)(23) xor ((not pi_in(1)(1)(23)) and pi_in(2)(2)(23));
 chi_out(0)(0)(24) <= pi_in(0)(0)(24) xor ((not pi_in(1)(1)(24)) and pi_in(2)(2)(24));
 chi_out(0)(0)(25) <= pi_in(0)(0)(25) xor ((not pi_in(1)(1)(25)) and pi_in(2)(2)(25));
 chi_out(0)(0)(26) <= pi_in(0)(0)(26) xor ((not pi_in(1)(1)(26)) and pi_in(2)(2)(26));
 chi_out(0)(0)(27) <= pi_in(0)(0)(27) xor ((not pi_in(1)(1)(27)) and pi_in(2)(2)(27));
 chi_out(0)(0)(28) <= pi_in(0)(0)(28) xor ((not pi_in(1)(1)(28)) and pi_in(2)(2)(28));
 chi_out(0)(0)(29) <= pi_in(0)(0)(29) xor ((not pi_in(1)(1)(29)) and pi_in(2)(2)(29));
 chi_out(0)(0)(30) <= pi_in(0)(0)(30) xor ((not pi_in(1)(1)(30)) and pi_in(2)(2)(30));
 chi_out(0)(0)(31) <= pi_in(0)(0)(31) xor ((not pi_in(1)(1)(31)) and pi_in(2)(2)(31));
 chi_out(0)(0)(32) <= pi_in(0)(0)(32) xor ((not pi_in(1)(1)(32)) and pi_in(2)(2)(32));
 chi_out(0)(0)(33) <= pi_in(0)(0)(33) xor ((not pi_in(1)(1)(33)) and pi_in(2)(2)(33));
 chi_out(0)(0)(34) <= pi_in(0)(0)(34) xor ((not pi_in(1)(1)(34)) and pi_in(2)(2)(34));
 chi_out(0)(0)(35) <= pi_in(0)(0)(35) xor ((not pi_in(1)(1)(35)) and pi_in(2)(2)(35));
 chi_out(0)(0)(36) <= pi_in(0)(0)(36) xor ((not pi_in(1)(1)(36)) and pi_in(2)(2)(36));
 chi_out(0)(0)(37) <= pi_in(0)(0)(37) xor ((not pi_in(1)(1)(37)) and pi_in(2)(2)(37));
 chi_out(0)(0)(38) <= pi_in(0)(0)(38) xor ((not pi_in(1)(1)(38)) and pi_in(2)(2)(38));
 chi_out(0)(0)(39) <= pi_in(0)(0)(39) xor ((not pi_in(1)(1)(39)) and pi_in(2)(2)(39));
 chi_out(0)(0)(40) <= pi_in(0)(0)(40) xor ((not pi_in(1)(1)(40)) and pi_in(2)(2)(40));
 chi_out(0)(0)(41) <= pi_in(0)(0)(41) xor ((not pi_in(1)(1)(41)) and pi_in(2)(2)(41));
 chi_out(0)(0)(42) <= pi_in(0)(0)(42) xor ((not pi_in(1)(1)(42)) and pi_in(2)(2)(42));
 chi_out(0)(0)(43) <= pi_in(0)(0)(43) xor ((not pi_in(1)(1)(43)) and pi_in(2)(2)(43));
 chi_out(0)(0)(44) <= pi_in(0)(0)(44) xor ((not pi_in(1)(1)(44)) and pi_in(2)(2)(44));
 chi_out(0)(0)(45) <= pi_in(0)(0)(45) xor ((not pi_in(1)(1)(45)) and pi_in(2)(2)(45));
 chi_out(0)(0)(46) <= pi_in(0)(0)(46) xor ((not pi_in(1)(1)(46)) and pi_in(2)(2)(46));
 chi_out(0)(0)(47) <= pi_in(0)(0)(47) xor ((not pi_in(1)(1)(47)) and pi_in(2)(2)(47));
 chi_out(0)(0)(48) <= pi_in(0)(0)(48) xor ((not pi_in(1)(1)(48)) and pi_in(2)(2)(48));
 chi_out(0)(0)(49) <= pi_in(0)(0)(49) xor ((not pi_in(1)(1)(49)) and pi_in(2)(2)(49));
 chi_out(0)(0)(50) <= pi_in(0)(0)(50) xor ((not pi_in(1)(1)(50)) and pi_in(2)(2)(50));
 chi_out(0)(0)(51) <= pi_in(0)(0)(51) xor ((not pi_in(1)(1)(51)) and pi_in(2)(2)(51));
 chi_out(0)(0)(52) <= pi_in(0)(0)(52) xor ((not pi_in(1)(1)(52)) and pi_in(2)(2)(52));
 chi_out(0)(0)(53) <= pi_in(0)(0)(53) xor ((not pi_in(1)(1)(53)) and pi_in(2)(2)(53));
 chi_out(0)(0)(54) <= pi_in(0)(0)(54) xor ((not pi_in(1)(1)(54)) and pi_in(2)(2)(54));
 chi_out(0)(0)(55) <= pi_in(0)(0)(55) xor ((not pi_in(1)(1)(55)) and pi_in(2)(2)(55));
 chi_out(0)(0)(56) <= pi_in(0)(0)(56) xor ((not pi_in(1)(1)(56)) and pi_in(2)(2)(56));
 chi_out(0)(0)(57) <= pi_in(0)(0)(57) xor ((not pi_in(1)(1)(57)) and pi_in(2)(2)(57));
 chi_out(0)(0)(58) <= pi_in(0)(0)(58) xor ((not pi_in(1)(1)(58)) and pi_in(2)(2)(58));
 chi_out(0)(0)(59) <= pi_in(0)(0)(59) xor ((not pi_in(1)(1)(59)) and pi_in(2)(2)(59));
 chi_out(0)(0)(60) <= pi_in(0)(0)(60) xor ((not pi_in(1)(1)(60)) and pi_in(2)(2)(60));
 chi_out(0)(0)(61) <= pi_in(0)(0)(61) xor ((not pi_in(1)(1)(61)) and pi_in(2)(2)(61));
 chi_out(0)(0)(62) <= pi_in(0)(0)(62) xor ((not pi_in(1)(1)(62)) and pi_in(2)(2)(62));
 chi_out(0)(0)(63) <= pi_in(0)(0)(63) xor ((not pi_in(1)(1)(63)) and pi_in(2)(2)(63));
 chi_out(0)(1)(0) <= pi_in(1)(1)(0) xor ((not pi_in(2)(2)(0)) and pi_in(3)(3)(0));
 chi_out(0)(1)(1) <= pi_in(1)(1)(1) xor ((not pi_in(2)(2)(1)) and pi_in(3)(3)(1));
 chi_out(0)(1)(2) <= pi_in(1)(1)(2) xor ((not pi_in(2)(2)(2)) and pi_in(3)(3)(2));
 chi_out(0)(1)(3) <= pi_in(1)(1)(3) xor ((not pi_in(2)(2)(3)) and pi_in(3)(3)(3));
 chi_out(0)(1)(4) <= pi_in(1)(1)(4) xor ((not pi_in(2)(2)(4)) and pi_in(3)(3)(4));
 chi_out(0)(1)(5) <= pi_in(1)(1)(5) xor ((not pi_in(2)(2)(5)) and pi_in(3)(3)(5));
 chi_out(0)(1)(6) <= pi_in(1)(1)(6) xor ((not pi_in(2)(2)(6)) and pi_in(3)(3)(6));
 chi_out(0)(1)(7) <= pi_in(1)(1)(7) xor ((not pi_in(2)(2)(7)) and pi_in(3)(3)(7));
 chi_out(0)(1)(8) <= pi_in(1)(1)(8) xor ((not pi_in(2)(2)(8)) and pi_in(3)(3)(8));
 chi_out(0)(1)(9) <= pi_in(1)(1)(9) xor ((not pi_in(2)(2)(9)) and pi_in(3)(3)(9));
 chi_out(0)(1)(10) <= pi_in(1)(1)(10) xor ((not pi_in(2)(2)(10)) and pi_in(3)(3)(10));
 chi_out(0)(1)(11) <= pi_in(1)(1)(11) xor ((not pi_in(2)(2)(11)) and pi_in(3)(3)(11));
 chi_out(0)(1)(12) <= pi_in(1)(1)(12) xor ((not pi_in(2)(2)(12)) and pi_in(3)(3)(12));
 chi_out(0)(1)(13) <= pi_in(1)(1)(13) xor ((not pi_in(2)(2)(13)) and pi_in(3)(3)(13));
 chi_out(0)(1)(14) <= pi_in(1)(1)(14) xor ((not pi_in(2)(2)(14)) and pi_in(3)(3)(14));
 chi_out(0)(1)(15) <= pi_in(1)(1)(15) xor ((not pi_in(2)(2)(15)) and pi_in(3)(3)(15));
 chi_out(0)(1)(16) <= pi_in(1)(1)(16) xor ((not pi_in(2)(2)(16)) and pi_in(3)(3)(16));
 chi_out(0)(1)(17) <= pi_in(1)(1)(17) xor ((not pi_in(2)(2)(17)) and pi_in(3)(3)(17));
 chi_out(0)(1)(18) <= pi_in(1)(1)(18) xor ((not pi_in(2)(2)(18)) and pi_in(3)(3)(18));
 chi_out(0)(1)(19) <= pi_in(1)(1)(19) xor ((not pi_in(2)(2)(19)) and pi_in(3)(3)(19));
 chi_out(0)(1)(20) <= pi_in(1)(1)(20) xor ((not pi_in(2)(2)(20)) and pi_in(3)(3)(20));
 chi_out(0)(1)(21) <= pi_in(1)(1)(21) xor ((not pi_in(2)(2)(21)) and pi_in(3)(3)(21));
 chi_out(0)(1)(22) <= pi_in(1)(1)(22) xor ((not pi_in(2)(2)(22)) and pi_in(3)(3)(22));
 chi_out(0)(1)(23) <= pi_in(1)(1)(23) xor ((not pi_in(2)(2)(23)) and pi_in(3)(3)(23));
 chi_out(0)(1)(24) <= pi_in(1)(1)(24) xor ((not pi_in(2)(2)(24)) and pi_in(3)(3)(24));
 chi_out(0)(1)(25) <= pi_in(1)(1)(25) xor ((not pi_in(2)(2)(25)) and pi_in(3)(3)(25));
 chi_out(0)(1)(26) <= pi_in(1)(1)(26) xor ((not pi_in(2)(2)(26)) and pi_in(3)(3)(26));
 chi_out(0)(1)(27) <= pi_in(1)(1)(27) xor ((not pi_in(2)(2)(27)) and pi_in(3)(3)(27));
 chi_out(0)(1)(28) <= pi_in(1)(1)(28) xor ((not pi_in(2)(2)(28)) and pi_in(3)(3)(28));
 chi_out(0)(1)(29) <= pi_in(1)(1)(29) xor ((not pi_in(2)(2)(29)) and pi_in(3)(3)(29));
 chi_out(0)(1)(30) <= pi_in(1)(1)(30) xor ((not pi_in(2)(2)(30)) and pi_in(3)(3)(30));
 chi_out(0)(1)(31) <= pi_in(1)(1)(31) xor ((not pi_in(2)(2)(31)) and pi_in(3)(3)(31));
 chi_out(0)(1)(32) <= pi_in(1)(1)(32) xor ((not pi_in(2)(2)(32)) and pi_in(3)(3)(32));
 chi_out(0)(1)(33) <= pi_in(1)(1)(33) xor ((not pi_in(2)(2)(33)) and pi_in(3)(3)(33));
 chi_out(0)(1)(34) <= pi_in(1)(1)(34) xor ((not pi_in(2)(2)(34)) and pi_in(3)(3)(34));
 chi_out(0)(1)(35) <= pi_in(1)(1)(35) xor ((not pi_in(2)(2)(35)) and pi_in(3)(3)(35));
 chi_out(0)(1)(36) <= pi_in(1)(1)(36) xor ((not pi_in(2)(2)(36)) and pi_in(3)(3)(36));
 chi_out(0)(1)(37) <= pi_in(1)(1)(37) xor ((not pi_in(2)(2)(37)) and pi_in(3)(3)(37));
 chi_out(0)(1)(38) <= pi_in(1)(1)(38) xor ((not pi_in(2)(2)(38)) and pi_in(3)(3)(38));
 chi_out(0)(1)(39) <= pi_in(1)(1)(39) xor ((not pi_in(2)(2)(39)) and pi_in(3)(3)(39));
 chi_out(0)(1)(40) <= pi_in(1)(1)(40) xor ((not pi_in(2)(2)(40)) and pi_in(3)(3)(40));
 chi_out(0)(1)(41) <= pi_in(1)(1)(41) xor ((not pi_in(2)(2)(41)) and pi_in(3)(3)(41));
 chi_out(0)(1)(42) <= pi_in(1)(1)(42) xor ((not pi_in(2)(2)(42)) and pi_in(3)(3)(42));
 chi_out(0)(1)(43) <= pi_in(1)(1)(43) xor ((not pi_in(2)(2)(43)) and pi_in(3)(3)(43));
 chi_out(0)(1)(44) <= pi_in(1)(1)(44) xor ((not pi_in(2)(2)(44)) and pi_in(3)(3)(44));
 chi_out(0)(1)(45) <= pi_in(1)(1)(45) xor ((not pi_in(2)(2)(45)) and pi_in(3)(3)(45));
 chi_out(0)(1)(46) <= pi_in(1)(1)(46) xor ((not pi_in(2)(2)(46)) and pi_in(3)(3)(46));
 chi_out(0)(1)(47) <= pi_in(1)(1)(47) xor ((not pi_in(2)(2)(47)) and pi_in(3)(3)(47));
 chi_out(0)(1)(48) <= pi_in(1)(1)(48) xor ((not pi_in(2)(2)(48)) and pi_in(3)(3)(48));
 chi_out(0)(1)(49) <= pi_in(1)(1)(49) xor ((not pi_in(2)(2)(49)) and pi_in(3)(3)(49));
 chi_out(0)(1)(50) <= pi_in(1)(1)(50) xor ((not pi_in(2)(2)(50)) and pi_in(3)(3)(50));
 chi_out(0)(1)(51) <= pi_in(1)(1)(51) xor ((not pi_in(2)(2)(51)) and pi_in(3)(3)(51));
 chi_out(0)(1)(52) <= pi_in(1)(1)(52) xor ((not pi_in(2)(2)(52)) and pi_in(3)(3)(52));
 chi_out(0)(1)(53) <= pi_in(1)(1)(53) xor ((not pi_in(2)(2)(53)) and pi_in(3)(3)(53));
 chi_out(0)(1)(54) <= pi_in(1)(1)(54) xor ((not pi_in(2)(2)(54)) and pi_in(3)(3)(54));
 chi_out(0)(1)(55) <= pi_in(1)(1)(55) xor ((not pi_in(2)(2)(55)) and pi_in(3)(3)(55));
 chi_out(0)(1)(56) <= pi_in(1)(1)(56) xor ((not pi_in(2)(2)(56)) and pi_in(3)(3)(56));
 chi_out(0)(1)(57) <= pi_in(1)(1)(57) xor ((not pi_in(2)(2)(57)) and pi_in(3)(3)(57));
 chi_out(0)(1)(58) <= pi_in(1)(1)(58) xor ((not pi_in(2)(2)(58)) and pi_in(3)(3)(58));
 chi_out(0)(1)(59) <= pi_in(1)(1)(59) xor ((not pi_in(2)(2)(59)) and pi_in(3)(3)(59));
 chi_out(0)(1)(60) <= pi_in(1)(1)(60) xor ((not pi_in(2)(2)(60)) and pi_in(3)(3)(60));
 chi_out(0)(1)(61) <= pi_in(1)(1)(61) xor ((not pi_in(2)(2)(61)) and pi_in(3)(3)(61));
 chi_out(0)(1)(62) <= pi_in(1)(1)(62) xor ((not pi_in(2)(2)(62)) and pi_in(3)(3)(62));
 chi_out(0)(1)(63) <= pi_in(1)(1)(63) xor ((not pi_in(2)(2)(63)) and pi_in(3)(3)(63));
 chi_out(0)(2)(0) <= pi_in(2)(2)(0) xor ((not pi_in(3)(3)(0)) and pi_in(4)(4)(0));
 chi_out(0)(2)(1) <= pi_in(2)(2)(1) xor ((not pi_in(3)(3)(1)) and pi_in(4)(4)(1));
 chi_out(0)(2)(2) <= pi_in(2)(2)(2) xor ((not pi_in(3)(3)(2)) and pi_in(4)(4)(2));
 chi_out(0)(2)(3) <= pi_in(2)(2)(3) xor ((not pi_in(3)(3)(3)) and pi_in(4)(4)(3));
 chi_out(0)(2)(4) <= pi_in(2)(2)(4) xor ((not pi_in(3)(3)(4)) and pi_in(4)(4)(4));
 chi_out(0)(2)(5) <= pi_in(2)(2)(5) xor ((not pi_in(3)(3)(5)) and pi_in(4)(4)(5));
 chi_out(0)(2)(6) <= pi_in(2)(2)(6) xor ((not pi_in(3)(3)(6)) and pi_in(4)(4)(6));
 chi_out(0)(2)(7) <= pi_in(2)(2)(7) xor ((not pi_in(3)(3)(7)) and pi_in(4)(4)(7));
 chi_out(0)(2)(8) <= pi_in(2)(2)(8) xor ((not pi_in(3)(3)(8)) and pi_in(4)(4)(8));
 chi_out(0)(2)(9) <= pi_in(2)(2)(9) xor ((not pi_in(3)(3)(9)) and pi_in(4)(4)(9));
 chi_out(0)(2)(10) <= pi_in(2)(2)(10) xor ((not pi_in(3)(3)(10)) and pi_in(4)(4)(10));
 chi_out(0)(2)(11) <= pi_in(2)(2)(11) xor ((not pi_in(3)(3)(11)) and pi_in(4)(4)(11));
 chi_out(0)(2)(12) <= pi_in(2)(2)(12) xor ((not pi_in(3)(3)(12)) and pi_in(4)(4)(12));
 chi_out(0)(2)(13) <= pi_in(2)(2)(13) xor ((not pi_in(3)(3)(13)) and pi_in(4)(4)(13));
 chi_out(0)(2)(14) <= pi_in(2)(2)(14) xor ((not pi_in(3)(3)(14)) and pi_in(4)(4)(14));
 chi_out(0)(2)(15) <= pi_in(2)(2)(15) xor ((not pi_in(3)(3)(15)) and pi_in(4)(4)(15));
 chi_out(0)(2)(16) <= pi_in(2)(2)(16) xor ((not pi_in(3)(3)(16)) and pi_in(4)(4)(16));
 chi_out(0)(2)(17) <= pi_in(2)(2)(17) xor ((not pi_in(3)(3)(17)) and pi_in(4)(4)(17));
 chi_out(0)(2)(18) <= pi_in(2)(2)(18) xor ((not pi_in(3)(3)(18)) and pi_in(4)(4)(18));
 chi_out(0)(2)(19) <= pi_in(2)(2)(19) xor ((not pi_in(3)(3)(19)) and pi_in(4)(4)(19));
 chi_out(0)(2)(20) <= pi_in(2)(2)(20) xor ((not pi_in(3)(3)(20)) and pi_in(4)(4)(20));
 chi_out(0)(2)(21) <= pi_in(2)(2)(21) xor ((not pi_in(3)(3)(21)) and pi_in(4)(4)(21));
 chi_out(0)(2)(22) <= pi_in(2)(2)(22) xor ((not pi_in(3)(3)(22)) and pi_in(4)(4)(22));
 chi_out(0)(2)(23) <= pi_in(2)(2)(23) xor ((not pi_in(3)(3)(23)) and pi_in(4)(4)(23));
 chi_out(0)(2)(24) <= pi_in(2)(2)(24) xor ((not pi_in(3)(3)(24)) and pi_in(4)(4)(24));
 chi_out(0)(2)(25) <= pi_in(2)(2)(25) xor ((not pi_in(3)(3)(25)) and pi_in(4)(4)(25));
 chi_out(0)(2)(26) <= pi_in(2)(2)(26) xor ((not pi_in(3)(3)(26)) and pi_in(4)(4)(26));
 chi_out(0)(2)(27) <= pi_in(2)(2)(27) xor ((not pi_in(3)(3)(27)) and pi_in(4)(4)(27));
 chi_out(0)(2)(28) <= pi_in(2)(2)(28) xor ((not pi_in(3)(3)(28)) and pi_in(4)(4)(28));
 chi_out(0)(2)(29) <= pi_in(2)(2)(29) xor ((not pi_in(3)(3)(29)) and pi_in(4)(4)(29));
 chi_out(0)(2)(30) <= pi_in(2)(2)(30) xor ((not pi_in(3)(3)(30)) and pi_in(4)(4)(30));
 chi_out(0)(2)(31) <= pi_in(2)(2)(31) xor ((not pi_in(3)(3)(31)) and pi_in(4)(4)(31));
 chi_out(0)(2)(32) <= pi_in(2)(2)(32) xor ((not pi_in(3)(3)(32)) and pi_in(4)(4)(32));
 chi_out(0)(2)(33) <= pi_in(2)(2)(33) xor ((not pi_in(3)(3)(33)) and pi_in(4)(4)(33));
 chi_out(0)(2)(34) <= pi_in(2)(2)(34) xor ((not pi_in(3)(3)(34)) and pi_in(4)(4)(34));
 chi_out(0)(2)(35) <= pi_in(2)(2)(35) xor ((not pi_in(3)(3)(35)) and pi_in(4)(4)(35));
 chi_out(0)(2)(36) <= pi_in(2)(2)(36) xor ((not pi_in(3)(3)(36)) and pi_in(4)(4)(36));
 chi_out(0)(2)(37) <= pi_in(2)(2)(37) xor ((not pi_in(3)(3)(37)) and pi_in(4)(4)(37));
 chi_out(0)(2)(38) <= pi_in(2)(2)(38) xor ((not pi_in(3)(3)(38)) and pi_in(4)(4)(38));
 chi_out(0)(2)(39) <= pi_in(2)(2)(39) xor ((not pi_in(3)(3)(39)) and pi_in(4)(4)(39));
 chi_out(0)(2)(40) <= pi_in(2)(2)(40) xor ((not pi_in(3)(3)(40)) and pi_in(4)(4)(40));
 chi_out(0)(2)(41) <= pi_in(2)(2)(41) xor ((not pi_in(3)(3)(41)) and pi_in(4)(4)(41));
 chi_out(0)(2)(42) <= pi_in(2)(2)(42) xor ((not pi_in(3)(3)(42)) and pi_in(4)(4)(42));
 chi_out(0)(2)(43) <= pi_in(2)(2)(43) xor ((not pi_in(3)(3)(43)) and pi_in(4)(4)(43));
 chi_out(0)(2)(44) <= pi_in(2)(2)(44) xor ((not pi_in(3)(3)(44)) and pi_in(4)(4)(44));
 chi_out(0)(2)(45) <= pi_in(2)(2)(45) xor ((not pi_in(3)(3)(45)) and pi_in(4)(4)(45));
 chi_out(0)(2)(46) <= pi_in(2)(2)(46) xor ((not pi_in(3)(3)(46)) and pi_in(4)(4)(46));
 chi_out(0)(2)(47) <= pi_in(2)(2)(47) xor ((not pi_in(3)(3)(47)) and pi_in(4)(4)(47));
 chi_out(0)(2)(48) <= pi_in(2)(2)(48) xor ((not pi_in(3)(3)(48)) and pi_in(4)(4)(48));
 chi_out(0)(2)(49) <= pi_in(2)(2)(49) xor ((not pi_in(3)(3)(49)) and pi_in(4)(4)(49));
 chi_out(0)(2)(50) <= pi_in(2)(2)(50) xor ((not pi_in(3)(3)(50)) and pi_in(4)(4)(50));
 chi_out(0)(2)(51) <= pi_in(2)(2)(51) xor ((not pi_in(3)(3)(51)) and pi_in(4)(4)(51));
 chi_out(0)(2)(52) <= pi_in(2)(2)(52) xor ((not pi_in(3)(3)(52)) and pi_in(4)(4)(52));
 chi_out(0)(2)(53) <= pi_in(2)(2)(53) xor ((not pi_in(3)(3)(53)) and pi_in(4)(4)(53));
 chi_out(0)(2)(54) <= pi_in(2)(2)(54) xor ((not pi_in(3)(3)(54)) and pi_in(4)(4)(54));
 chi_out(0)(2)(55) <= pi_in(2)(2)(55) xor ((not pi_in(3)(3)(55)) and pi_in(4)(4)(55));
 chi_out(0)(2)(56) <= pi_in(2)(2)(56) xor ((not pi_in(3)(3)(56)) and pi_in(4)(4)(56));
 chi_out(0)(2)(57) <= pi_in(2)(2)(57) xor ((not pi_in(3)(3)(57)) and pi_in(4)(4)(57));
 chi_out(0)(2)(58) <= pi_in(2)(2)(58) xor ((not pi_in(3)(3)(58)) and pi_in(4)(4)(58));
 chi_out(0)(2)(59) <= pi_in(2)(2)(59) xor ((not pi_in(3)(3)(59)) and pi_in(4)(4)(59));
 chi_out(0)(2)(60) <= pi_in(2)(2)(60) xor ((not pi_in(3)(3)(60)) and pi_in(4)(4)(60));
 chi_out(0)(2)(61) <= pi_in(2)(2)(61) xor ((not pi_in(3)(3)(61)) and pi_in(4)(4)(61));
 chi_out(0)(2)(62) <= pi_in(2)(2)(62) xor ((not pi_in(3)(3)(62)) and pi_in(4)(4)(62));
 chi_out(0)(2)(63) <= pi_in(2)(2)(63) xor ((not pi_in(3)(3)(63)) and pi_in(4)(4)(63));
 chi_out(1)(0)(0) <= pi_in(0)(3)(0) xor ((not pi_in(1)(4)(0)) and pi_in(2)(0)(0));
 chi_out(1)(0)(1) <= pi_in(0)(3)(1) xor ((not pi_in(1)(4)(1)) and pi_in(2)(0)(1));
 chi_out(1)(0)(2) <= pi_in(0)(3)(2) xor ((not pi_in(1)(4)(2)) and pi_in(2)(0)(2));
 chi_out(1)(0)(3) <= pi_in(0)(3)(3) xor ((not pi_in(1)(4)(3)) and pi_in(2)(0)(3));
 chi_out(1)(0)(4) <= pi_in(0)(3)(4) xor ((not pi_in(1)(4)(4)) and pi_in(2)(0)(4));
 chi_out(1)(0)(5) <= pi_in(0)(3)(5) xor ((not pi_in(1)(4)(5)) and pi_in(2)(0)(5));
 chi_out(1)(0)(6) <= pi_in(0)(3)(6) xor ((not pi_in(1)(4)(6)) and pi_in(2)(0)(6));
 chi_out(1)(0)(7) <= pi_in(0)(3)(7) xor ((not pi_in(1)(4)(7)) and pi_in(2)(0)(7));
 chi_out(1)(0)(8) <= pi_in(0)(3)(8) xor ((not pi_in(1)(4)(8)) and pi_in(2)(0)(8));
 chi_out(1)(0)(9) <= pi_in(0)(3)(9) xor ((not pi_in(1)(4)(9)) and pi_in(2)(0)(9));
 chi_out(1)(0)(10) <= pi_in(0)(3)(10) xor ((not pi_in(1)(4)(10)) and pi_in(2)(0)(10));
 chi_out(1)(0)(11) <= pi_in(0)(3)(11) xor ((not pi_in(1)(4)(11)) and pi_in(2)(0)(11));
 chi_out(1)(0)(12) <= pi_in(0)(3)(12) xor ((not pi_in(1)(4)(12)) and pi_in(2)(0)(12));
 chi_out(1)(0)(13) <= pi_in(0)(3)(13) xor ((not pi_in(1)(4)(13)) and pi_in(2)(0)(13));
 chi_out(1)(0)(14) <= pi_in(0)(3)(14) xor ((not pi_in(1)(4)(14)) and pi_in(2)(0)(14));
 chi_out(1)(0)(15) <= pi_in(0)(3)(15) xor ((not pi_in(1)(4)(15)) and pi_in(2)(0)(15));
 chi_out(1)(0)(16) <= pi_in(0)(3)(16) xor ((not pi_in(1)(4)(16)) and pi_in(2)(0)(16));
 chi_out(1)(0)(17) <= pi_in(0)(3)(17) xor ((not pi_in(1)(4)(17)) and pi_in(2)(0)(17));
 chi_out(1)(0)(18) <= pi_in(0)(3)(18) xor ((not pi_in(1)(4)(18)) and pi_in(2)(0)(18));
 chi_out(1)(0)(19) <= pi_in(0)(3)(19) xor ((not pi_in(1)(4)(19)) and pi_in(2)(0)(19));
 chi_out(1)(0)(20) <= pi_in(0)(3)(20) xor ((not pi_in(1)(4)(20)) and pi_in(2)(0)(20));
 chi_out(1)(0)(21) <= pi_in(0)(3)(21) xor ((not pi_in(1)(4)(21)) and pi_in(2)(0)(21));
 chi_out(1)(0)(22) <= pi_in(0)(3)(22) xor ((not pi_in(1)(4)(22)) and pi_in(2)(0)(22));
 chi_out(1)(0)(23) <= pi_in(0)(3)(23) xor ((not pi_in(1)(4)(23)) and pi_in(2)(0)(23));
 chi_out(1)(0)(24) <= pi_in(0)(3)(24) xor ((not pi_in(1)(4)(24)) and pi_in(2)(0)(24));
 chi_out(1)(0)(25) <= pi_in(0)(3)(25) xor ((not pi_in(1)(4)(25)) and pi_in(2)(0)(25));
 chi_out(1)(0)(26) <= pi_in(0)(3)(26) xor ((not pi_in(1)(4)(26)) and pi_in(2)(0)(26));
 chi_out(1)(0)(27) <= pi_in(0)(3)(27) xor ((not pi_in(1)(4)(27)) and pi_in(2)(0)(27));
 chi_out(1)(0)(28) <= pi_in(0)(3)(28) xor ((not pi_in(1)(4)(28)) and pi_in(2)(0)(28));
 chi_out(1)(0)(29) <= pi_in(0)(3)(29) xor ((not pi_in(1)(4)(29)) and pi_in(2)(0)(29));
 chi_out(1)(0)(30) <= pi_in(0)(3)(30) xor ((not pi_in(1)(4)(30)) and pi_in(2)(0)(30));
 chi_out(1)(0)(31) <= pi_in(0)(3)(31) xor ((not pi_in(1)(4)(31)) and pi_in(2)(0)(31));
 chi_out(1)(0)(32) <= pi_in(0)(3)(32) xor ((not pi_in(1)(4)(32)) and pi_in(2)(0)(32));
 chi_out(1)(0)(33) <= pi_in(0)(3)(33) xor ((not pi_in(1)(4)(33)) and pi_in(2)(0)(33));
 chi_out(1)(0)(34) <= pi_in(0)(3)(34) xor ((not pi_in(1)(4)(34)) and pi_in(2)(0)(34));
 chi_out(1)(0)(35) <= pi_in(0)(3)(35) xor ((not pi_in(1)(4)(35)) and pi_in(2)(0)(35));
 chi_out(1)(0)(36) <= pi_in(0)(3)(36) xor ((not pi_in(1)(4)(36)) and pi_in(2)(0)(36));
 chi_out(1)(0)(37) <= pi_in(0)(3)(37) xor ((not pi_in(1)(4)(37)) and pi_in(2)(0)(37));
 chi_out(1)(0)(38) <= pi_in(0)(3)(38) xor ((not pi_in(1)(4)(38)) and pi_in(2)(0)(38));
 chi_out(1)(0)(39) <= pi_in(0)(3)(39) xor ((not pi_in(1)(4)(39)) and pi_in(2)(0)(39));
 chi_out(1)(0)(40) <= pi_in(0)(3)(40) xor ((not pi_in(1)(4)(40)) and pi_in(2)(0)(40));
 chi_out(1)(0)(41) <= pi_in(0)(3)(41) xor ((not pi_in(1)(4)(41)) and pi_in(2)(0)(41));
 chi_out(1)(0)(42) <= pi_in(0)(3)(42) xor ((not pi_in(1)(4)(42)) and pi_in(2)(0)(42));
 chi_out(1)(0)(43) <= pi_in(0)(3)(43) xor ((not pi_in(1)(4)(43)) and pi_in(2)(0)(43));
 chi_out(1)(0)(44) <= pi_in(0)(3)(44) xor ((not pi_in(1)(4)(44)) and pi_in(2)(0)(44));
 chi_out(1)(0)(45) <= pi_in(0)(3)(45) xor ((not pi_in(1)(4)(45)) and pi_in(2)(0)(45));
 chi_out(1)(0)(46) <= pi_in(0)(3)(46) xor ((not pi_in(1)(4)(46)) and pi_in(2)(0)(46));
 chi_out(1)(0)(47) <= pi_in(0)(3)(47) xor ((not pi_in(1)(4)(47)) and pi_in(2)(0)(47));
 chi_out(1)(0)(48) <= pi_in(0)(3)(48) xor ((not pi_in(1)(4)(48)) and pi_in(2)(0)(48));
 chi_out(1)(0)(49) <= pi_in(0)(3)(49) xor ((not pi_in(1)(4)(49)) and pi_in(2)(0)(49));
 chi_out(1)(0)(50) <= pi_in(0)(3)(50) xor ((not pi_in(1)(4)(50)) and pi_in(2)(0)(50));
 chi_out(1)(0)(51) <= pi_in(0)(3)(51) xor ((not pi_in(1)(4)(51)) and pi_in(2)(0)(51));
 chi_out(1)(0)(52) <= pi_in(0)(3)(52) xor ((not pi_in(1)(4)(52)) and pi_in(2)(0)(52));
 chi_out(1)(0)(53) <= pi_in(0)(3)(53) xor ((not pi_in(1)(4)(53)) and pi_in(2)(0)(53));
 chi_out(1)(0)(54) <= pi_in(0)(3)(54) xor ((not pi_in(1)(4)(54)) and pi_in(2)(0)(54));
 chi_out(1)(0)(55) <= pi_in(0)(3)(55) xor ((not pi_in(1)(4)(55)) and pi_in(2)(0)(55));
 chi_out(1)(0)(56) <= pi_in(0)(3)(56) xor ((not pi_in(1)(4)(56)) and pi_in(2)(0)(56));
 chi_out(1)(0)(57) <= pi_in(0)(3)(57) xor ((not pi_in(1)(4)(57)) and pi_in(2)(0)(57));
 chi_out(1)(0)(58) <= pi_in(0)(3)(58) xor ((not pi_in(1)(4)(58)) and pi_in(2)(0)(58));
 chi_out(1)(0)(59) <= pi_in(0)(3)(59) xor ((not pi_in(1)(4)(59)) and pi_in(2)(0)(59));
 chi_out(1)(0)(60) <= pi_in(0)(3)(60) xor ((not pi_in(1)(4)(60)) and pi_in(2)(0)(60));
 chi_out(1)(0)(61) <= pi_in(0)(3)(61) xor ((not pi_in(1)(4)(61)) and pi_in(2)(0)(61));
 chi_out(1)(0)(62) <= pi_in(0)(3)(62) xor ((not pi_in(1)(4)(62)) and pi_in(2)(0)(62));
 chi_out(1)(0)(63) <= pi_in(0)(3)(63) xor ((not pi_in(1)(4)(63)) and pi_in(2)(0)(63));
 chi_out(1)(1)(0) <= pi_in(1)(4)(0) xor ((not pi_in(2)(0)(0)) and pi_in(3)(1)(0));
 chi_out(1)(1)(1) <= pi_in(1)(4)(1) xor ((not pi_in(2)(0)(1)) and pi_in(3)(1)(1));
 chi_out(1)(1)(2) <= pi_in(1)(4)(2) xor ((not pi_in(2)(0)(2)) and pi_in(3)(1)(2));
 chi_out(1)(1)(3) <= pi_in(1)(4)(3) xor ((not pi_in(2)(0)(3)) and pi_in(3)(1)(3));
 chi_out(1)(1)(4) <= pi_in(1)(4)(4) xor ((not pi_in(2)(0)(4)) and pi_in(3)(1)(4));
 chi_out(1)(1)(5) <= pi_in(1)(4)(5) xor ((not pi_in(2)(0)(5)) and pi_in(3)(1)(5));
 chi_out(1)(1)(6) <= pi_in(1)(4)(6) xor ((not pi_in(2)(0)(6)) and pi_in(3)(1)(6));
 chi_out(1)(1)(7) <= pi_in(1)(4)(7) xor ((not pi_in(2)(0)(7)) and pi_in(3)(1)(7));
 chi_out(1)(1)(8) <= pi_in(1)(4)(8) xor ((not pi_in(2)(0)(8)) and pi_in(3)(1)(8));
 chi_out(1)(1)(9) <= pi_in(1)(4)(9) xor ((not pi_in(2)(0)(9)) and pi_in(3)(1)(9));
 chi_out(1)(1)(10) <= pi_in(1)(4)(10) xor ((not pi_in(2)(0)(10)) and pi_in(3)(1)(10));
 chi_out(1)(1)(11) <= pi_in(1)(4)(11) xor ((not pi_in(2)(0)(11)) and pi_in(3)(1)(11));
 chi_out(1)(1)(12) <= pi_in(1)(4)(12) xor ((not pi_in(2)(0)(12)) and pi_in(3)(1)(12));
 chi_out(1)(1)(13) <= pi_in(1)(4)(13) xor ((not pi_in(2)(0)(13)) and pi_in(3)(1)(13));
 chi_out(1)(1)(14) <= pi_in(1)(4)(14) xor ((not pi_in(2)(0)(14)) and pi_in(3)(1)(14));
 chi_out(1)(1)(15) <= pi_in(1)(4)(15) xor ((not pi_in(2)(0)(15)) and pi_in(3)(1)(15));
 chi_out(1)(1)(16) <= pi_in(1)(4)(16) xor ((not pi_in(2)(0)(16)) and pi_in(3)(1)(16));
 chi_out(1)(1)(17) <= pi_in(1)(4)(17) xor ((not pi_in(2)(0)(17)) and pi_in(3)(1)(17));
 chi_out(1)(1)(18) <= pi_in(1)(4)(18) xor ((not pi_in(2)(0)(18)) and pi_in(3)(1)(18));
 chi_out(1)(1)(19) <= pi_in(1)(4)(19) xor ((not pi_in(2)(0)(19)) and pi_in(3)(1)(19));
 chi_out(1)(1)(20) <= pi_in(1)(4)(20) xor ((not pi_in(2)(0)(20)) and pi_in(3)(1)(20));
 chi_out(1)(1)(21) <= pi_in(1)(4)(21) xor ((not pi_in(2)(0)(21)) and pi_in(3)(1)(21));
 chi_out(1)(1)(22) <= pi_in(1)(4)(22) xor ((not pi_in(2)(0)(22)) and pi_in(3)(1)(22));
 chi_out(1)(1)(23) <= pi_in(1)(4)(23) xor ((not pi_in(2)(0)(23)) and pi_in(3)(1)(23));
 chi_out(1)(1)(24) <= pi_in(1)(4)(24) xor ((not pi_in(2)(0)(24)) and pi_in(3)(1)(24));
 chi_out(1)(1)(25) <= pi_in(1)(4)(25) xor ((not pi_in(2)(0)(25)) and pi_in(3)(1)(25));
 chi_out(1)(1)(26) <= pi_in(1)(4)(26) xor ((not pi_in(2)(0)(26)) and pi_in(3)(1)(26));
 chi_out(1)(1)(27) <= pi_in(1)(4)(27) xor ((not pi_in(2)(0)(27)) and pi_in(3)(1)(27));
 chi_out(1)(1)(28) <= pi_in(1)(4)(28) xor ((not pi_in(2)(0)(28)) and pi_in(3)(1)(28));
 chi_out(1)(1)(29) <= pi_in(1)(4)(29) xor ((not pi_in(2)(0)(29)) and pi_in(3)(1)(29));
 chi_out(1)(1)(30) <= pi_in(1)(4)(30) xor ((not pi_in(2)(0)(30)) and pi_in(3)(1)(30));
 chi_out(1)(1)(31) <= pi_in(1)(4)(31) xor ((not pi_in(2)(0)(31)) and pi_in(3)(1)(31));
 chi_out(1)(1)(32) <= pi_in(1)(4)(32) xor ((not pi_in(2)(0)(32)) and pi_in(3)(1)(32));
 chi_out(1)(1)(33) <= pi_in(1)(4)(33) xor ((not pi_in(2)(0)(33)) and pi_in(3)(1)(33));
 chi_out(1)(1)(34) <= pi_in(1)(4)(34) xor ((not pi_in(2)(0)(34)) and pi_in(3)(1)(34));
 chi_out(1)(1)(35) <= pi_in(1)(4)(35) xor ((not pi_in(2)(0)(35)) and pi_in(3)(1)(35));
 chi_out(1)(1)(36) <= pi_in(1)(4)(36) xor ((not pi_in(2)(0)(36)) and pi_in(3)(1)(36));
 chi_out(1)(1)(37) <= pi_in(1)(4)(37) xor ((not pi_in(2)(0)(37)) and pi_in(3)(1)(37));
 chi_out(1)(1)(38) <= pi_in(1)(4)(38) xor ((not pi_in(2)(0)(38)) and pi_in(3)(1)(38));
 chi_out(1)(1)(39) <= pi_in(1)(4)(39) xor ((not pi_in(2)(0)(39)) and pi_in(3)(1)(39));
 chi_out(1)(1)(40) <= pi_in(1)(4)(40) xor ((not pi_in(2)(0)(40)) and pi_in(3)(1)(40));
 chi_out(1)(1)(41) <= pi_in(1)(4)(41) xor ((not pi_in(2)(0)(41)) and pi_in(3)(1)(41));
 chi_out(1)(1)(42) <= pi_in(1)(4)(42) xor ((not pi_in(2)(0)(42)) and pi_in(3)(1)(42));
 chi_out(1)(1)(43) <= pi_in(1)(4)(43) xor ((not pi_in(2)(0)(43)) and pi_in(3)(1)(43));
 chi_out(1)(1)(44) <= pi_in(1)(4)(44) xor ((not pi_in(2)(0)(44)) and pi_in(3)(1)(44));
 chi_out(1)(1)(45) <= pi_in(1)(4)(45) xor ((not pi_in(2)(0)(45)) and pi_in(3)(1)(45));
 chi_out(1)(1)(46) <= pi_in(1)(4)(46) xor ((not pi_in(2)(0)(46)) and pi_in(3)(1)(46));
 chi_out(1)(1)(47) <= pi_in(1)(4)(47) xor ((not pi_in(2)(0)(47)) and pi_in(3)(1)(47));
 chi_out(1)(1)(48) <= pi_in(1)(4)(48) xor ((not pi_in(2)(0)(48)) and pi_in(3)(1)(48));
 chi_out(1)(1)(49) <= pi_in(1)(4)(49) xor ((not pi_in(2)(0)(49)) and pi_in(3)(1)(49));
 chi_out(1)(1)(50) <= pi_in(1)(4)(50) xor ((not pi_in(2)(0)(50)) and pi_in(3)(1)(50));
 chi_out(1)(1)(51) <= pi_in(1)(4)(51) xor ((not pi_in(2)(0)(51)) and pi_in(3)(1)(51));
 chi_out(1)(1)(52) <= pi_in(1)(4)(52) xor ((not pi_in(2)(0)(52)) and pi_in(3)(1)(52));
 chi_out(1)(1)(53) <= pi_in(1)(4)(53) xor ((not pi_in(2)(0)(53)) and pi_in(3)(1)(53));
 chi_out(1)(1)(54) <= pi_in(1)(4)(54) xor ((not pi_in(2)(0)(54)) and pi_in(3)(1)(54));
 chi_out(1)(1)(55) <= pi_in(1)(4)(55) xor ((not pi_in(2)(0)(55)) and pi_in(3)(1)(55));
 chi_out(1)(1)(56) <= pi_in(1)(4)(56) xor ((not pi_in(2)(0)(56)) and pi_in(3)(1)(56));
 chi_out(1)(1)(57) <= pi_in(1)(4)(57) xor ((not pi_in(2)(0)(57)) and pi_in(3)(1)(57));
 chi_out(1)(1)(58) <= pi_in(1)(4)(58) xor ((not pi_in(2)(0)(58)) and pi_in(3)(1)(58));
 chi_out(1)(1)(59) <= pi_in(1)(4)(59) xor ((not pi_in(2)(0)(59)) and pi_in(3)(1)(59));
 chi_out(1)(1)(60) <= pi_in(1)(4)(60) xor ((not pi_in(2)(0)(60)) and pi_in(3)(1)(60));
 chi_out(1)(1)(61) <= pi_in(1)(4)(61) xor ((not pi_in(2)(0)(61)) and pi_in(3)(1)(61));
 chi_out(1)(1)(62) <= pi_in(1)(4)(62) xor ((not pi_in(2)(0)(62)) and pi_in(3)(1)(62));
 chi_out(1)(1)(63) <= pi_in(1)(4)(63) xor ((not pi_in(2)(0)(63)) and pi_in(3)(1)(63));
 chi_out(1)(2)(0) <= pi_in(2)(0)(0) xor ((not pi_in(3)(1)(0)) and pi_in(4)(2)(0));
 chi_out(1)(2)(1) <= pi_in(2)(0)(1) xor ((not pi_in(3)(1)(1)) and pi_in(4)(2)(1));
 chi_out(1)(2)(2) <= pi_in(2)(0)(2) xor ((not pi_in(3)(1)(2)) and pi_in(4)(2)(2));
 chi_out(1)(2)(3) <= pi_in(2)(0)(3) xor ((not pi_in(3)(1)(3)) and pi_in(4)(2)(3));
 chi_out(1)(2)(4) <= pi_in(2)(0)(4) xor ((not pi_in(3)(1)(4)) and pi_in(4)(2)(4));
 chi_out(1)(2)(5) <= pi_in(2)(0)(5) xor ((not pi_in(3)(1)(5)) and pi_in(4)(2)(5));
 chi_out(1)(2)(6) <= pi_in(2)(0)(6) xor ((not pi_in(3)(1)(6)) and pi_in(4)(2)(6));
 chi_out(1)(2)(7) <= pi_in(2)(0)(7) xor ((not pi_in(3)(1)(7)) and pi_in(4)(2)(7));
 chi_out(1)(2)(8) <= pi_in(2)(0)(8) xor ((not pi_in(3)(1)(8)) and pi_in(4)(2)(8));
 chi_out(1)(2)(9) <= pi_in(2)(0)(9) xor ((not pi_in(3)(1)(9)) and pi_in(4)(2)(9));
 chi_out(1)(2)(10) <= pi_in(2)(0)(10) xor ((not pi_in(3)(1)(10)) and pi_in(4)(2)(10));
 chi_out(1)(2)(11) <= pi_in(2)(0)(11) xor ((not pi_in(3)(1)(11)) and pi_in(4)(2)(11));
 chi_out(1)(2)(12) <= pi_in(2)(0)(12) xor ((not pi_in(3)(1)(12)) and pi_in(4)(2)(12));
 chi_out(1)(2)(13) <= pi_in(2)(0)(13) xor ((not pi_in(3)(1)(13)) and pi_in(4)(2)(13));
 chi_out(1)(2)(14) <= pi_in(2)(0)(14) xor ((not pi_in(3)(1)(14)) and pi_in(4)(2)(14));
 chi_out(1)(2)(15) <= pi_in(2)(0)(15) xor ((not pi_in(3)(1)(15)) and pi_in(4)(2)(15));
 chi_out(1)(2)(16) <= pi_in(2)(0)(16) xor ((not pi_in(3)(1)(16)) and pi_in(4)(2)(16));
 chi_out(1)(2)(17) <= pi_in(2)(0)(17) xor ((not pi_in(3)(1)(17)) and pi_in(4)(2)(17));
 chi_out(1)(2)(18) <= pi_in(2)(0)(18) xor ((not pi_in(3)(1)(18)) and pi_in(4)(2)(18));
 chi_out(1)(2)(19) <= pi_in(2)(0)(19) xor ((not pi_in(3)(1)(19)) and pi_in(4)(2)(19));
 chi_out(1)(2)(20) <= pi_in(2)(0)(20) xor ((not pi_in(3)(1)(20)) and pi_in(4)(2)(20));
 chi_out(1)(2)(21) <= pi_in(2)(0)(21) xor ((not pi_in(3)(1)(21)) and pi_in(4)(2)(21));
 chi_out(1)(2)(22) <= pi_in(2)(0)(22) xor ((not pi_in(3)(1)(22)) and pi_in(4)(2)(22));
 chi_out(1)(2)(23) <= pi_in(2)(0)(23) xor ((not pi_in(3)(1)(23)) and pi_in(4)(2)(23));
 chi_out(1)(2)(24) <= pi_in(2)(0)(24) xor ((not pi_in(3)(1)(24)) and pi_in(4)(2)(24));
 chi_out(1)(2)(25) <= pi_in(2)(0)(25) xor ((not pi_in(3)(1)(25)) and pi_in(4)(2)(25));
 chi_out(1)(2)(26) <= pi_in(2)(0)(26) xor ((not pi_in(3)(1)(26)) and pi_in(4)(2)(26));
 chi_out(1)(2)(27) <= pi_in(2)(0)(27) xor ((not pi_in(3)(1)(27)) and pi_in(4)(2)(27));
 chi_out(1)(2)(28) <= pi_in(2)(0)(28) xor ((not pi_in(3)(1)(28)) and pi_in(4)(2)(28));
 chi_out(1)(2)(29) <= pi_in(2)(0)(29) xor ((not pi_in(3)(1)(29)) and pi_in(4)(2)(29));
 chi_out(1)(2)(30) <= pi_in(2)(0)(30) xor ((not pi_in(3)(1)(30)) and pi_in(4)(2)(30));
 chi_out(1)(2)(31) <= pi_in(2)(0)(31) xor ((not pi_in(3)(1)(31)) and pi_in(4)(2)(31));
 chi_out(1)(2)(32) <= pi_in(2)(0)(32) xor ((not pi_in(3)(1)(32)) and pi_in(4)(2)(32));
 chi_out(1)(2)(33) <= pi_in(2)(0)(33) xor ((not pi_in(3)(1)(33)) and pi_in(4)(2)(33));
 chi_out(1)(2)(34) <= pi_in(2)(0)(34) xor ((not pi_in(3)(1)(34)) and pi_in(4)(2)(34));
 chi_out(1)(2)(35) <= pi_in(2)(0)(35) xor ((not pi_in(3)(1)(35)) and pi_in(4)(2)(35));
 chi_out(1)(2)(36) <= pi_in(2)(0)(36) xor ((not pi_in(3)(1)(36)) and pi_in(4)(2)(36));
 chi_out(1)(2)(37) <= pi_in(2)(0)(37) xor ((not pi_in(3)(1)(37)) and pi_in(4)(2)(37));
 chi_out(1)(2)(38) <= pi_in(2)(0)(38) xor ((not pi_in(3)(1)(38)) and pi_in(4)(2)(38));
 chi_out(1)(2)(39) <= pi_in(2)(0)(39) xor ((not pi_in(3)(1)(39)) and pi_in(4)(2)(39));
 chi_out(1)(2)(40) <= pi_in(2)(0)(40) xor ((not pi_in(3)(1)(40)) and pi_in(4)(2)(40));
 chi_out(1)(2)(41) <= pi_in(2)(0)(41) xor ((not pi_in(3)(1)(41)) and pi_in(4)(2)(41));
 chi_out(1)(2)(42) <= pi_in(2)(0)(42) xor ((not pi_in(3)(1)(42)) and pi_in(4)(2)(42));
 chi_out(1)(2)(43) <= pi_in(2)(0)(43) xor ((not pi_in(3)(1)(43)) and pi_in(4)(2)(43));
 chi_out(1)(2)(44) <= pi_in(2)(0)(44) xor ((not pi_in(3)(1)(44)) and pi_in(4)(2)(44));
 chi_out(1)(2)(45) <= pi_in(2)(0)(45) xor ((not pi_in(3)(1)(45)) and pi_in(4)(2)(45));
 chi_out(1)(2)(46) <= pi_in(2)(0)(46) xor ((not pi_in(3)(1)(46)) and pi_in(4)(2)(46));
 chi_out(1)(2)(47) <= pi_in(2)(0)(47) xor ((not pi_in(3)(1)(47)) and pi_in(4)(2)(47));
 chi_out(1)(2)(48) <= pi_in(2)(0)(48) xor ((not pi_in(3)(1)(48)) and pi_in(4)(2)(48));
 chi_out(1)(2)(49) <= pi_in(2)(0)(49) xor ((not pi_in(3)(1)(49)) and pi_in(4)(2)(49));
 chi_out(1)(2)(50) <= pi_in(2)(0)(50) xor ((not pi_in(3)(1)(50)) and pi_in(4)(2)(50));
 chi_out(1)(2)(51) <= pi_in(2)(0)(51) xor ((not pi_in(3)(1)(51)) and pi_in(4)(2)(51));
 chi_out(1)(2)(52) <= pi_in(2)(0)(52) xor ((not pi_in(3)(1)(52)) and pi_in(4)(2)(52));
 chi_out(1)(2)(53) <= pi_in(2)(0)(53) xor ((not pi_in(3)(1)(53)) and pi_in(4)(2)(53));
 chi_out(1)(2)(54) <= pi_in(2)(0)(54) xor ((not pi_in(3)(1)(54)) and pi_in(4)(2)(54));
 chi_out(1)(2)(55) <= pi_in(2)(0)(55) xor ((not pi_in(3)(1)(55)) and pi_in(4)(2)(55));
 chi_out(1)(2)(56) <= pi_in(2)(0)(56) xor ((not pi_in(3)(1)(56)) and pi_in(4)(2)(56));
 chi_out(1)(2)(57) <= pi_in(2)(0)(57) xor ((not pi_in(3)(1)(57)) and pi_in(4)(2)(57));
 chi_out(1)(2)(58) <= pi_in(2)(0)(58) xor ((not pi_in(3)(1)(58)) and pi_in(4)(2)(58));
 chi_out(1)(2)(59) <= pi_in(2)(0)(59) xor ((not pi_in(3)(1)(59)) and pi_in(4)(2)(59));
 chi_out(1)(2)(60) <= pi_in(2)(0)(60) xor ((not pi_in(3)(1)(60)) and pi_in(4)(2)(60));
 chi_out(1)(2)(61) <= pi_in(2)(0)(61) xor ((not pi_in(3)(1)(61)) and pi_in(4)(2)(61));
 chi_out(1)(2)(62) <= pi_in(2)(0)(62) xor ((not pi_in(3)(1)(62)) and pi_in(4)(2)(62));
 chi_out(1)(2)(63) <= pi_in(2)(0)(63) xor ((not pi_in(3)(1)(63)) and pi_in(4)(2)(63));
 chi_out(2)(0)(0) <= pi_in(0)(1)(0) xor ((not pi_in(1)(2)(0)) and pi_in(2)(3)(0));
 chi_out(2)(0)(1) <= pi_in(0)(1)(1) xor ((not pi_in(1)(2)(1)) and pi_in(2)(3)(1));
 chi_out(2)(0)(2) <= pi_in(0)(1)(2) xor ((not pi_in(1)(2)(2)) and pi_in(2)(3)(2));
 chi_out(2)(0)(3) <= pi_in(0)(1)(3) xor ((not pi_in(1)(2)(3)) and pi_in(2)(3)(3));
 chi_out(2)(0)(4) <= pi_in(0)(1)(4) xor ((not pi_in(1)(2)(4)) and pi_in(2)(3)(4));
 chi_out(2)(0)(5) <= pi_in(0)(1)(5) xor ((not pi_in(1)(2)(5)) and pi_in(2)(3)(5));
 chi_out(2)(0)(6) <= pi_in(0)(1)(6) xor ((not pi_in(1)(2)(6)) and pi_in(2)(3)(6));
 chi_out(2)(0)(7) <= pi_in(0)(1)(7) xor ((not pi_in(1)(2)(7)) and pi_in(2)(3)(7));
 chi_out(2)(0)(8) <= pi_in(0)(1)(8) xor ((not pi_in(1)(2)(8)) and pi_in(2)(3)(8));
 chi_out(2)(0)(9) <= pi_in(0)(1)(9) xor ((not pi_in(1)(2)(9)) and pi_in(2)(3)(9));
 chi_out(2)(0)(10) <= pi_in(0)(1)(10) xor ((not pi_in(1)(2)(10)) and pi_in(2)(3)(10));
 chi_out(2)(0)(11) <= pi_in(0)(1)(11) xor ((not pi_in(1)(2)(11)) and pi_in(2)(3)(11));
 chi_out(2)(0)(12) <= pi_in(0)(1)(12) xor ((not pi_in(1)(2)(12)) and pi_in(2)(3)(12));
 chi_out(2)(0)(13) <= pi_in(0)(1)(13) xor ((not pi_in(1)(2)(13)) and pi_in(2)(3)(13));
 chi_out(2)(0)(14) <= pi_in(0)(1)(14) xor ((not pi_in(1)(2)(14)) and pi_in(2)(3)(14));
 chi_out(2)(0)(15) <= pi_in(0)(1)(15) xor ((not pi_in(1)(2)(15)) and pi_in(2)(3)(15));
 chi_out(2)(0)(16) <= pi_in(0)(1)(16) xor ((not pi_in(1)(2)(16)) and pi_in(2)(3)(16));
 chi_out(2)(0)(17) <= pi_in(0)(1)(17) xor ((not pi_in(1)(2)(17)) and pi_in(2)(3)(17));
 chi_out(2)(0)(18) <= pi_in(0)(1)(18) xor ((not pi_in(1)(2)(18)) and pi_in(2)(3)(18));
 chi_out(2)(0)(19) <= pi_in(0)(1)(19) xor ((not pi_in(1)(2)(19)) and pi_in(2)(3)(19));
 chi_out(2)(0)(20) <= pi_in(0)(1)(20) xor ((not pi_in(1)(2)(20)) and pi_in(2)(3)(20));
 chi_out(2)(0)(21) <= pi_in(0)(1)(21) xor ((not pi_in(1)(2)(21)) and pi_in(2)(3)(21));
 chi_out(2)(0)(22) <= pi_in(0)(1)(22) xor ((not pi_in(1)(2)(22)) and pi_in(2)(3)(22));
 chi_out(2)(0)(23) <= pi_in(0)(1)(23) xor ((not pi_in(1)(2)(23)) and pi_in(2)(3)(23));
 chi_out(2)(0)(24) <= pi_in(0)(1)(24) xor ((not pi_in(1)(2)(24)) and pi_in(2)(3)(24));
 chi_out(2)(0)(25) <= pi_in(0)(1)(25) xor ((not pi_in(1)(2)(25)) and pi_in(2)(3)(25));
 chi_out(2)(0)(26) <= pi_in(0)(1)(26) xor ((not pi_in(1)(2)(26)) and pi_in(2)(3)(26));
 chi_out(2)(0)(27) <= pi_in(0)(1)(27) xor ((not pi_in(1)(2)(27)) and pi_in(2)(3)(27));
 chi_out(2)(0)(28) <= pi_in(0)(1)(28) xor ((not pi_in(1)(2)(28)) and pi_in(2)(3)(28));
 chi_out(2)(0)(29) <= pi_in(0)(1)(29) xor ((not pi_in(1)(2)(29)) and pi_in(2)(3)(29));
 chi_out(2)(0)(30) <= pi_in(0)(1)(30) xor ((not pi_in(1)(2)(30)) and pi_in(2)(3)(30));
 chi_out(2)(0)(31) <= pi_in(0)(1)(31) xor ((not pi_in(1)(2)(31)) and pi_in(2)(3)(31));
 chi_out(2)(0)(32) <= pi_in(0)(1)(32) xor ((not pi_in(1)(2)(32)) and pi_in(2)(3)(32));
 chi_out(2)(0)(33) <= pi_in(0)(1)(33) xor ((not pi_in(1)(2)(33)) and pi_in(2)(3)(33));
 chi_out(2)(0)(34) <= pi_in(0)(1)(34) xor ((not pi_in(1)(2)(34)) and pi_in(2)(3)(34));
 chi_out(2)(0)(35) <= pi_in(0)(1)(35) xor ((not pi_in(1)(2)(35)) and pi_in(2)(3)(35));
 chi_out(2)(0)(36) <= pi_in(0)(1)(36) xor ((not pi_in(1)(2)(36)) and pi_in(2)(3)(36));
 chi_out(2)(0)(37) <= pi_in(0)(1)(37) xor ((not pi_in(1)(2)(37)) and pi_in(2)(3)(37));
 chi_out(2)(0)(38) <= pi_in(0)(1)(38) xor ((not pi_in(1)(2)(38)) and pi_in(2)(3)(38));
 chi_out(2)(0)(39) <= pi_in(0)(1)(39) xor ((not pi_in(1)(2)(39)) and pi_in(2)(3)(39));
 chi_out(2)(0)(40) <= pi_in(0)(1)(40) xor ((not pi_in(1)(2)(40)) and pi_in(2)(3)(40));
 chi_out(2)(0)(41) <= pi_in(0)(1)(41) xor ((not pi_in(1)(2)(41)) and pi_in(2)(3)(41));
 chi_out(2)(0)(42) <= pi_in(0)(1)(42) xor ((not pi_in(1)(2)(42)) and pi_in(2)(3)(42));
 chi_out(2)(0)(43) <= pi_in(0)(1)(43) xor ((not pi_in(1)(2)(43)) and pi_in(2)(3)(43));
 chi_out(2)(0)(44) <= pi_in(0)(1)(44) xor ((not pi_in(1)(2)(44)) and pi_in(2)(3)(44));
 chi_out(2)(0)(45) <= pi_in(0)(1)(45) xor ((not pi_in(1)(2)(45)) and pi_in(2)(3)(45));
 chi_out(2)(0)(46) <= pi_in(0)(1)(46) xor ((not pi_in(1)(2)(46)) and pi_in(2)(3)(46));
 chi_out(2)(0)(47) <= pi_in(0)(1)(47) xor ((not pi_in(1)(2)(47)) and pi_in(2)(3)(47));
 chi_out(2)(0)(48) <= pi_in(0)(1)(48) xor ((not pi_in(1)(2)(48)) and pi_in(2)(3)(48));
 chi_out(2)(0)(49) <= pi_in(0)(1)(49) xor ((not pi_in(1)(2)(49)) and pi_in(2)(3)(49));
 chi_out(2)(0)(50) <= pi_in(0)(1)(50) xor ((not pi_in(1)(2)(50)) and pi_in(2)(3)(50));
 chi_out(2)(0)(51) <= pi_in(0)(1)(51) xor ((not pi_in(1)(2)(51)) and pi_in(2)(3)(51));
 chi_out(2)(0)(52) <= pi_in(0)(1)(52) xor ((not pi_in(1)(2)(52)) and pi_in(2)(3)(52));
 chi_out(2)(0)(53) <= pi_in(0)(1)(53) xor ((not pi_in(1)(2)(53)) and pi_in(2)(3)(53));
 chi_out(2)(0)(54) <= pi_in(0)(1)(54) xor ((not pi_in(1)(2)(54)) and pi_in(2)(3)(54));
 chi_out(2)(0)(55) <= pi_in(0)(1)(55) xor ((not pi_in(1)(2)(55)) and pi_in(2)(3)(55));
 chi_out(2)(0)(56) <= pi_in(0)(1)(56) xor ((not pi_in(1)(2)(56)) and pi_in(2)(3)(56));
 chi_out(2)(0)(57) <= pi_in(0)(1)(57) xor ((not pi_in(1)(2)(57)) and pi_in(2)(3)(57));
 chi_out(2)(0)(58) <= pi_in(0)(1)(58) xor ((not pi_in(1)(2)(58)) and pi_in(2)(3)(58));
 chi_out(2)(0)(59) <= pi_in(0)(1)(59) xor ((not pi_in(1)(2)(59)) and pi_in(2)(3)(59));
 chi_out(2)(0)(60) <= pi_in(0)(1)(60) xor ((not pi_in(1)(2)(60)) and pi_in(2)(3)(60));
 chi_out(2)(0)(61) <= pi_in(0)(1)(61) xor ((not pi_in(1)(2)(61)) and pi_in(2)(3)(61));
 chi_out(2)(0)(62) <= pi_in(0)(1)(62) xor ((not pi_in(1)(2)(62)) and pi_in(2)(3)(62));
 chi_out(2)(0)(63) <= pi_in(0)(1)(63) xor ((not pi_in(1)(2)(63)) and pi_in(2)(3)(63));
 chi_out(2)(1)(0) <= pi_in(1)(2)(0) xor ((not pi_in(2)(3)(0)) and pi_in(3)(4)(0));
 chi_out(2)(1)(1) <= pi_in(1)(2)(1) xor ((not pi_in(2)(3)(1)) and pi_in(3)(4)(1));
 chi_out(2)(1)(2) <= pi_in(1)(2)(2) xor ((not pi_in(2)(3)(2)) and pi_in(3)(4)(2));
 chi_out(2)(1)(3) <= pi_in(1)(2)(3) xor ((not pi_in(2)(3)(3)) and pi_in(3)(4)(3));
 chi_out(2)(1)(4) <= pi_in(1)(2)(4) xor ((not pi_in(2)(3)(4)) and pi_in(3)(4)(4));
 chi_out(2)(1)(5) <= pi_in(1)(2)(5) xor ((not pi_in(2)(3)(5)) and pi_in(3)(4)(5));
 chi_out(2)(1)(6) <= pi_in(1)(2)(6) xor ((not pi_in(2)(3)(6)) and pi_in(3)(4)(6));
 chi_out(2)(1)(7) <= pi_in(1)(2)(7) xor ((not pi_in(2)(3)(7)) and pi_in(3)(4)(7));
 chi_out(2)(1)(8) <= pi_in(1)(2)(8) xor ((not pi_in(2)(3)(8)) and pi_in(3)(4)(8));
 chi_out(2)(1)(9) <= pi_in(1)(2)(9) xor ((not pi_in(2)(3)(9)) and pi_in(3)(4)(9));
 chi_out(2)(1)(10) <= pi_in(1)(2)(10) xor ((not pi_in(2)(3)(10)) and pi_in(3)(4)(10));
 chi_out(2)(1)(11) <= pi_in(1)(2)(11) xor ((not pi_in(2)(3)(11)) and pi_in(3)(4)(11));
 chi_out(2)(1)(12) <= pi_in(1)(2)(12) xor ((not pi_in(2)(3)(12)) and pi_in(3)(4)(12));
 chi_out(2)(1)(13) <= pi_in(1)(2)(13) xor ((not pi_in(2)(3)(13)) and pi_in(3)(4)(13));
 chi_out(2)(1)(14) <= pi_in(1)(2)(14) xor ((not pi_in(2)(3)(14)) and pi_in(3)(4)(14));
 chi_out(2)(1)(15) <= pi_in(1)(2)(15) xor ((not pi_in(2)(3)(15)) and pi_in(3)(4)(15));
 chi_out(2)(1)(16) <= pi_in(1)(2)(16) xor ((not pi_in(2)(3)(16)) and pi_in(3)(4)(16));
 chi_out(2)(1)(17) <= pi_in(1)(2)(17) xor ((not pi_in(2)(3)(17)) and pi_in(3)(4)(17));
 chi_out(2)(1)(18) <= pi_in(1)(2)(18) xor ((not pi_in(2)(3)(18)) and pi_in(3)(4)(18));
 chi_out(2)(1)(19) <= pi_in(1)(2)(19) xor ((not pi_in(2)(3)(19)) and pi_in(3)(4)(19));
 chi_out(2)(1)(20) <= pi_in(1)(2)(20) xor ((not pi_in(2)(3)(20)) and pi_in(3)(4)(20));
 chi_out(2)(1)(21) <= pi_in(1)(2)(21) xor ((not pi_in(2)(3)(21)) and pi_in(3)(4)(21));
 chi_out(2)(1)(22) <= pi_in(1)(2)(22) xor ((not pi_in(2)(3)(22)) and pi_in(3)(4)(22));
 chi_out(2)(1)(23) <= pi_in(1)(2)(23) xor ((not pi_in(2)(3)(23)) and pi_in(3)(4)(23));
 chi_out(2)(1)(24) <= pi_in(1)(2)(24) xor ((not pi_in(2)(3)(24)) and pi_in(3)(4)(24));
 chi_out(2)(1)(25) <= pi_in(1)(2)(25) xor ((not pi_in(2)(3)(25)) and pi_in(3)(4)(25));
 chi_out(2)(1)(26) <= pi_in(1)(2)(26) xor ((not pi_in(2)(3)(26)) and pi_in(3)(4)(26));
 chi_out(2)(1)(27) <= pi_in(1)(2)(27) xor ((not pi_in(2)(3)(27)) and pi_in(3)(4)(27));
 chi_out(2)(1)(28) <= pi_in(1)(2)(28) xor ((not pi_in(2)(3)(28)) and pi_in(3)(4)(28));
 chi_out(2)(1)(29) <= pi_in(1)(2)(29) xor ((not pi_in(2)(3)(29)) and pi_in(3)(4)(29));
 chi_out(2)(1)(30) <= pi_in(1)(2)(30) xor ((not pi_in(2)(3)(30)) and pi_in(3)(4)(30));
 chi_out(2)(1)(31) <= pi_in(1)(2)(31) xor ((not pi_in(2)(3)(31)) and pi_in(3)(4)(31));
 chi_out(2)(1)(32) <= pi_in(1)(2)(32) xor ((not pi_in(2)(3)(32)) and pi_in(3)(4)(32));
 chi_out(2)(1)(33) <= pi_in(1)(2)(33) xor ((not pi_in(2)(3)(33)) and pi_in(3)(4)(33));
 chi_out(2)(1)(34) <= pi_in(1)(2)(34) xor ((not pi_in(2)(3)(34)) and pi_in(3)(4)(34));
 chi_out(2)(1)(35) <= pi_in(1)(2)(35) xor ((not pi_in(2)(3)(35)) and pi_in(3)(4)(35));
 chi_out(2)(1)(36) <= pi_in(1)(2)(36) xor ((not pi_in(2)(3)(36)) and pi_in(3)(4)(36));
 chi_out(2)(1)(37) <= pi_in(1)(2)(37) xor ((not pi_in(2)(3)(37)) and pi_in(3)(4)(37));
 chi_out(2)(1)(38) <= pi_in(1)(2)(38) xor ((not pi_in(2)(3)(38)) and pi_in(3)(4)(38));
 chi_out(2)(1)(39) <= pi_in(1)(2)(39) xor ((not pi_in(2)(3)(39)) and pi_in(3)(4)(39));
 chi_out(2)(1)(40) <= pi_in(1)(2)(40) xor ((not pi_in(2)(3)(40)) and pi_in(3)(4)(40));
 chi_out(2)(1)(41) <= pi_in(1)(2)(41) xor ((not pi_in(2)(3)(41)) and pi_in(3)(4)(41));
 chi_out(2)(1)(42) <= pi_in(1)(2)(42) xor ((not pi_in(2)(3)(42)) and pi_in(3)(4)(42));
 chi_out(2)(1)(43) <= pi_in(1)(2)(43) xor ((not pi_in(2)(3)(43)) and pi_in(3)(4)(43));
 chi_out(2)(1)(44) <= pi_in(1)(2)(44) xor ((not pi_in(2)(3)(44)) and pi_in(3)(4)(44));
 chi_out(2)(1)(45) <= pi_in(1)(2)(45) xor ((not pi_in(2)(3)(45)) and pi_in(3)(4)(45));
 chi_out(2)(1)(46) <= pi_in(1)(2)(46) xor ((not pi_in(2)(3)(46)) and pi_in(3)(4)(46));
 chi_out(2)(1)(47) <= pi_in(1)(2)(47) xor ((not pi_in(2)(3)(47)) and pi_in(3)(4)(47));
 chi_out(2)(1)(48) <= pi_in(1)(2)(48) xor ((not pi_in(2)(3)(48)) and pi_in(3)(4)(48));
 chi_out(2)(1)(49) <= pi_in(1)(2)(49) xor ((not pi_in(2)(3)(49)) and pi_in(3)(4)(49));
 chi_out(2)(1)(50) <= pi_in(1)(2)(50) xor ((not pi_in(2)(3)(50)) and pi_in(3)(4)(50));
 chi_out(2)(1)(51) <= pi_in(1)(2)(51) xor ((not pi_in(2)(3)(51)) and pi_in(3)(4)(51));
 chi_out(2)(1)(52) <= pi_in(1)(2)(52) xor ((not pi_in(2)(3)(52)) and pi_in(3)(4)(52));
 chi_out(2)(1)(53) <= pi_in(1)(2)(53) xor ((not pi_in(2)(3)(53)) and pi_in(3)(4)(53));
 chi_out(2)(1)(54) <= pi_in(1)(2)(54) xor ((not pi_in(2)(3)(54)) and pi_in(3)(4)(54));
 chi_out(2)(1)(55) <= pi_in(1)(2)(55) xor ((not pi_in(2)(3)(55)) and pi_in(3)(4)(55));
 chi_out(2)(1)(56) <= pi_in(1)(2)(56) xor ((not pi_in(2)(3)(56)) and pi_in(3)(4)(56));
 chi_out(2)(1)(57) <= pi_in(1)(2)(57) xor ((not pi_in(2)(3)(57)) and pi_in(3)(4)(57));
 chi_out(2)(1)(58) <= pi_in(1)(2)(58) xor ((not pi_in(2)(3)(58)) and pi_in(3)(4)(58));
 chi_out(2)(1)(59) <= pi_in(1)(2)(59) xor ((not pi_in(2)(3)(59)) and pi_in(3)(4)(59));
 chi_out(2)(1)(60) <= pi_in(1)(2)(60) xor ((not pi_in(2)(3)(60)) and pi_in(3)(4)(60));
 chi_out(2)(1)(61) <= pi_in(1)(2)(61) xor ((not pi_in(2)(3)(61)) and pi_in(3)(4)(61));
 chi_out(2)(1)(62) <= pi_in(1)(2)(62) xor ((not pi_in(2)(3)(62)) and pi_in(3)(4)(62));
 chi_out(2)(1)(63) <= pi_in(1)(2)(63) xor ((not pi_in(2)(3)(63)) and pi_in(3)(4)(63));
 chi_out(2)(2)(0) <= pi_in(2)(3)(0) xor ((not pi_in(3)(4)(0)) and pi_in(4)(0)(0));
 chi_out(2)(2)(1) <= pi_in(2)(3)(1) xor ((not pi_in(3)(4)(1)) and pi_in(4)(0)(1));
 chi_out(2)(2)(2) <= pi_in(2)(3)(2) xor ((not pi_in(3)(4)(2)) and pi_in(4)(0)(2));
 chi_out(2)(2)(3) <= pi_in(2)(3)(3) xor ((not pi_in(3)(4)(3)) and pi_in(4)(0)(3));
 chi_out(2)(2)(4) <= pi_in(2)(3)(4) xor ((not pi_in(3)(4)(4)) and pi_in(4)(0)(4));
 chi_out(2)(2)(5) <= pi_in(2)(3)(5) xor ((not pi_in(3)(4)(5)) and pi_in(4)(0)(5));
 chi_out(2)(2)(6) <= pi_in(2)(3)(6) xor ((not pi_in(3)(4)(6)) and pi_in(4)(0)(6));
 chi_out(2)(2)(7) <= pi_in(2)(3)(7) xor ((not pi_in(3)(4)(7)) and pi_in(4)(0)(7));
 chi_out(2)(2)(8) <= pi_in(2)(3)(8) xor ((not pi_in(3)(4)(8)) and pi_in(4)(0)(8));
 chi_out(2)(2)(9) <= pi_in(2)(3)(9) xor ((not pi_in(3)(4)(9)) and pi_in(4)(0)(9));
 chi_out(2)(2)(10) <= pi_in(2)(3)(10) xor ((not pi_in(3)(4)(10)) and pi_in(4)(0)(10));
 chi_out(2)(2)(11) <= pi_in(2)(3)(11) xor ((not pi_in(3)(4)(11)) and pi_in(4)(0)(11));
 chi_out(2)(2)(12) <= pi_in(2)(3)(12) xor ((not pi_in(3)(4)(12)) and pi_in(4)(0)(12));
 chi_out(2)(2)(13) <= pi_in(2)(3)(13) xor ((not pi_in(3)(4)(13)) and pi_in(4)(0)(13));
 chi_out(2)(2)(14) <= pi_in(2)(3)(14) xor ((not pi_in(3)(4)(14)) and pi_in(4)(0)(14));
 chi_out(2)(2)(15) <= pi_in(2)(3)(15) xor ((not pi_in(3)(4)(15)) and pi_in(4)(0)(15));
 chi_out(2)(2)(16) <= pi_in(2)(3)(16) xor ((not pi_in(3)(4)(16)) and pi_in(4)(0)(16));
 chi_out(2)(2)(17) <= pi_in(2)(3)(17) xor ((not pi_in(3)(4)(17)) and pi_in(4)(0)(17));
 chi_out(2)(2)(18) <= pi_in(2)(3)(18) xor ((not pi_in(3)(4)(18)) and pi_in(4)(0)(18));
 chi_out(2)(2)(19) <= pi_in(2)(3)(19) xor ((not pi_in(3)(4)(19)) and pi_in(4)(0)(19));
 chi_out(2)(2)(20) <= pi_in(2)(3)(20) xor ((not pi_in(3)(4)(20)) and pi_in(4)(0)(20));
 chi_out(2)(2)(21) <= pi_in(2)(3)(21) xor ((not pi_in(3)(4)(21)) and pi_in(4)(0)(21));
 chi_out(2)(2)(22) <= pi_in(2)(3)(22) xor ((not pi_in(3)(4)(22)) and pi_in(4)(0)(22));
 chi_out(2)(2)(23) <= pi_in(2)(3)(23) xor ((not pi_in(3)(4)(23)) and pi_in(4)(0)(23));
 chi_out(2)(2)(24) <= pi_in(2)(3)(24) xor ((not pi_in(3)(4)(24)) and pi_in(4)(0)(24));
 chi_out(2)(2)(25) <= pi_in(2)(3)(25) xor ((not pi_in(3)(4)(25)) and pi_in(4)(0)(25));
 chi_out(2)(2)(26) <= pi_in(2)(3)(26) xor ((not pi_in(3)(4)(26)) and pi_in(4)(0)(26));
 chi_out(2)(2)(27) <= pi_in(2)(3)(27) xor ((not pi_in(3)(4)(27)) and pi_in(4)(0)(27));
 chi_out(2)(2)(28) <= pi_in(2)(3)(28) xor ((not pi_in(3)(4)(28)) and pi_in(4)(0)(28));
 chi_out(2)(2)(29) <= pi_in(2)(3)(29) xor ((not pi_in(3)(4)(29)) and pi_in(4)(0)(29));
 chi_out(2)(2)(30) <= pi_in(2)(3)(30) xor ((not pi_in(3)(4)(30)) and pi_in(4)(0)(30));
 chi_out(2)(2)(31) <= pi_in(2)(3)(31) xor ((not pi_in(3)(4)(31)) and pi_in(4)(0)(31));
 chi_out(2)(2)(32) <= pi_in(2)(3)(32) xor ((not pi_in(3)(4)(32)) and pi_in(4)(0)(32));
 chi_out(2)(2)(33) <= pi_in(2)(3)(33) xor ((not pi_in(3)(4)(33)) and pi_in(4)(0)(33));
 chi_out(2)(2)(34) <= pi_in(2)(3)(34) xor ((not pi_in(3)(4)(34)) and pi_in(4)(0)(34));
 chi_out(2)(2)(35) <= pi_in(2)(3)(35) xor ((not pi_in(3)(4)(35)) and pi_in(4)(0)(35));
 chi_out(2)(2)(36) <= pi_in(2)(3)(36) xor ((not pi_in(3)(4)(36)) and pi_in(4)(0)(36));
 chi_out(2)(2)(37) <= pi_in(2)(3)(37) xor ((not pi_in(3)(4)(37)) and pi_in(4)(0)(37));
 chi_out(2)(2)(38) <= pi_in(2)(3)(38) xor ((not pi_in(3)(4)(38)) and pi_in(4)(0)(38));
 chi_out(2)(2)(39) <= pi_in(2)(3)(39) xor ((not pi_in(3)(4)(39)) and pi_in(4)(0)(39));
 chi_out(2)(2)(40) <= pi_in(2)(3)(40) xor ((not pi_in(3)(4)(40)) and pi_in(4)(0)(40));
 chi_out(2)(2)(41) <= pi_in(2)(3)(41) xor ((not pi_in(3)(4)(41)) and pi_in(4)(0)(41));
 chi_out(2)(2)(42) <= pi_in(2)(3)(42) xor ((not pi_in(3)(4)(42)) and pi_in(4)(0)(42));
 chi_out(2)(2)(43) <= pi_in(2)(3)(43) xor ((not pi_in(3)(4)(43)) and pi_in(4)(0)(43));
 chi_out(2)(2)(44) <= pi_in(2)(3)(44) xor ((not pi_in(3)(4)(44)) and pi_in(4)(0)(44));
 chi_out(2)(2)(45) <= pi_in(2)(3)(45) xor ((not pi_in(3)(4)(45)) and pi_in(4)(0)(45));
 chi_out(2)(2)(46) <= pi_in(2)(3)(46) xor ((not pi_in(3)(4)(46)) and pi_in(4)(0)(46));
 chi_out(2)(2)(47) <= pi_in(2)(3)(47) xor ((not pi_in(3)(4)(47)) and pi_in(4)(0)(47));
 chi_out(2)(2)(48) <= pi_in(2)(3)(48) xor ((not pi_in(3)(4)(48)) and pi_in(4)(0)(48));
 chi_out(2)(2)(49) <= pi_in(2)(3)(49) xor ((not pi_in(3)(4)(49)) and pi_in(4)(0)(49));
 chi_out(2)(2)(50) <= pi_in(2)(3)(50) xor ((not pi_in(3)(4)(50)) and pi_in(4)(0)(50));
 chi_out(2)(2)(51) <= pi_in(2)(3)(51) xor ((not pi_in(3)(4)(51)) and pi_in(4)(0)(51));
 chi_out(2)(2)(52) <= pi_in(2)(3)(52) xor ((not pi_in(3)(4)(52)) and pi_in(4)(0)(52));
 chi_out(2)(2)(53) <= pi_in(2)(3)(53) xor ((not pi_in(3)(4)(53)) and pi_in(4)(0)(53));
 chi_out(2)(2)(54) <= pi_in(2)(3)(54) xor ((not pi_in(3)(4)(54)) and pi_in(4)(0)(54));
 chi_out(2)(2)(55) <= pi_in(2)(3)(55) xor ((not pi_in(3)(4)(55)) and pi_in(4)(0)(55));
 chi_out(2)(2)(56) <= pi_in(2)(3)(56) xor ((not pi_in(3)(4)(56)) and pi_in(4)(0)(56));
 chi_out(2)(2)(57) <= pi_in(2)(3)(57) xor ((not pi_in(3)(4)(57)) and pi_in(4)(0)(57));
 chi_out(2)(2)(58) <= pi_in(2)(3)(58) xor ((not pi_in(3)(4)(58)) and pi_in(4)(0)(58));
 chi_out(2)(2)(59) <= pi_in(2)(3)(59) xor ((not pi_in(3)(4)(59)) and pi_in(4)(0)(59));
 chi_out(2)(2)(60) <= pi_in(2)(3)(60) xor ((not pi_in(3)(4)(60)) and pi_in(4)(0)(60));
 chi_out(2)(2)(61) <= pi_in(2)(3)(61) xor ((not pi_in(3)(4)(61)) and pi_in(4)(0)(61));
 chi_out(2)(2)(62) <= pi_in(2)(3)(62) xor ((not pi_in(3)(4)(62)) and pi_in(4)(0)(62));
 chi_out(2)(2)(63) <= pi_in(2)(3)(63) xor ((not pi_in(3)(4)(63)) and pi_in(4)(0)(63));
 chi_out(3)(0)(0) <= pi_in(0)(4)(0) xor ((not pi_in(1)(0)(0)) and pi_in(2)(1)(0));
 chi_out(3)(0)(1) <= pi_in(0)(4)(1) xor ((not pi_in(1)(0)(1)) and pi_in(2)(1)(1));
 chi_out(3)(0)(2) <= pi_in(0)(4)(2) xor ((not pi_in(1)(0)(2)) and pi_in(2)(1)(2));
 chi_out(3)(0)(3) <= pi_in(0)(4)(3) xor ((not pi_in(1)(0)(3)) and pi_in(2)(1)(3));
 chi_out(3)(0)(4) <= pi_in(0)(4)(4) xor ((not pi_in(1)(0)(4)) and pi_in(2)(1)(4));
 chi_out(3)(0)(5) <= pi_in(0)(4)(5) xor ((not pi_in(1)(0)(5)) and pi_in(2)(1)(5));
 chi_out(3)(0)(6) <= pi_in(0)(4)(6) xor ((not pi_in(1)(0)(6)) and pi_in(2)(1)(6));
 chi_out(3)(0)(7) <= pi_in(0)(4)(7) xor ((not pi_in(1)(0)(7)) and pi_in(2)(1)(7));
 chi_out(3)(0)(8) <= pi_in(0)(4)(8) xor ((not pi_in(1)(0)(8)) and pi_in(2)(1)(8));
 chi_out(3)(0)(9) <= pi_in(0)(4)(9) xor ((not pi_in(1)(0)(9)) and pi_in(2)(1)(9));
 chi_out(3)(0)(10) <= pi_in(0)(4)(10) xor ((not pi_in(1)(0)(10)) and pi_in(2)(1)(10));
 chi_out(3)(0)(11) <= pi_in(0)(4)(11) xor ((not pi_in(1)(0)(11)) and pi_in(2)(1)(11));
 chi_out(3)(0)(12) <= pi_in(0)(4)(12) xor ((not pi_in(1)(0)(12)) and pi_in(2)(1)(12));
 chi_out(3)(0)(13) <= pi_in(0)(4)(13) xor ((not pi_in(1)(0)(13)) and pi_in(2)(1)(13));
 chi_out(3)(0)(14) <= pi_in(0)(4)(14) xor ((not pi_in(1)(0)(14)) and pi_in(2)(1)(14));
 chi_out(3)(0)(15) <= pi_in(0)(4)(15) xor ((not pi_in(1)(0)(15)) and pi_in(2)(1)(15));
 chi_out(3)(0)(16) <= pi_in(0)(4)(16) xor ((not pi_in(1)(0)(16)) and pi_in(2)(1)(16));
 chi_out(3)(0)(17) <= pi_in(0)(4)(17) xor ((not pi_in(1)(0)(17)) and pi_in(2)(1)(17));
 chi_out(3)(0)(18) <= pi_in(0)(4)(18) xor ((not pi_in(1)(0)(18)) and pi_in(2)(1)(18));
 chi_out(3)(0)(19) <= pi_in(0)(4)(19) xor ((not pi_in(1)(0)(19)) and pi_in(2)(1)(19));
 chi_out(3)(0)(20) <= pi_in(0)(4)(20) xor ((not pi_in(1)(0)(20)) and pi_in(2)(1)(20));
 chi_out(3)(0)(21) <= pi_in(0)(4)(21) xor ((not pi_in(1)(0)(21)) and pi_in(2)(1)(21));
 chi_out(3)(0)(22) <= pi_in(0)(4)(22) xor ((not pi_in(1)(0)(22)) and pi_in(2)(1)(22));
 chi_out(3)(0)(23) <= pi_in(0)(4)(23) xor ((not pi_in(1)(0)(23)) and pi_in(2)(1)(23));
 chi_out(3)(0)(24) <= pi_in(0)(4)(24) xor ((not pi_in(1)(0)(24)) and pi_in(2)(1)(24));
 chi_out(3)(0)(25) <= pi_in(0)(4)(25) xor ((not pi_in(1)(0)(25)) and pi_in(2)(1)(25));
 chi_out(3)(0)(26) <= pi_in(0)(4)(26) xor ((not pi_in(1)(0)(26)) and pi_in(2)(1)(26));
 chi_out(3)(0)(27) <= pi_in(0)(4)(27) xor ((not pi_in(1)(0)(27)) and pi_in(2)(1)(27));
 chi_out(3)(0)(28) <= pi_in(0)(4)(28) xor ((not pi_in(1)(0)(28)) and pi_in(2)(1)(28));
 chi_out(3)(0)(29) <= pi_in(0)(4)(29) xor ((not pi_in(1)(0)(29)) and pi_in(2)(1)(29));
 chi_out(3)(0)(30) <= pi_in(0)(4)(30) xor ((not pi_in(1)(0)(30)) and pi_in(2)(1)(30));
 chi_out(3)(0)(31) <= pi_in(0)(4)(31) xor ((not pi_in(1)(0)(31)) and pi_in(2)(1)(31));
 chi_out(3)(0)(32) <= pi_in(0)(4)(32) xor ((not pi_in(1)(0)(32)) and pi_in(2)(1)(32));
 chi_out(3)(0)(33) <= pi_in(0)(4)(33) xor ((not pi_in(1)(0)(33)) and pi_in(2)(1)(33));
 chi_out(3)(0)(34) <= pi_in(0)(4)(34) xor ((not pi_in(1)(0)(34)) and pi_in(2)(1)(34));
 chi_out(3)(0)(35) <= pi_in(0)(4)(35) xor ((not pi_in(1)(0)(35)) and pi_in(2)(1)(35));
 chi_out(3)(0)(36) <= pi_in(0)(4)(36) xor ((not pi_in(1)(0)(36)) and pi_in(2)(1)(36));
 chi_out(3)(0)(37) <= pi_in(0)(4)(37) xor ((not pi_in(1)(0)(37)) and pi_in(2)(1)(37));
 chi_out(3)(0)(38) <= pi_in(0)(4)(38) xor ((not pi_in(1)(0)(38)) and pi_in(2)(1)(38));
 chi_out(3)(0)(39) <= pi_in(0)(4)(39) xor ((not pi_in(1)(0)(39)) and pi_in(2)(1)(39));
 chi_out(3)(0)(40) <= pi_in(0)(4)(40) xor ((not pi_in(1)(0)(40)) and pi_in(2)(1)(40));
 chi_out(3)(0)(41) <= pi_in(0)(4)(41) xor ((not pi_in(1)(0)(41)) and pi_in(2)(1)(41));
 chi_out(3)(0)(42) <= pi_in(0)(4)(42) xor ((not pi_in(1)(0)(42)) and pi_in(2)(1)(42));
 chi_out(3)(0)(43) <= pi_in(0)(4)(43) xor ((not pi_in(1)(0)(43)) and pi_in(2)(1)(43));
 chi_out(3)(0)(44) <= pi_in(0)(4)(44) xor ((not pi_in(1)(0)(44)) and pi_in(2)(1)(44));
 chi_out(3)(0)(45) <= pi_in(0)(4)(45) xor ((not pi_in(1)(0)(45)) and pi_in(2)(1)(45));
 chi_out(3)(0)(46) <= pi_in(0)(4)(46) xor ((not pi_in(1)(0)(46)) and pi_in(2)(1)(46));
 chi_out(3)(0)(47) <= pi_in(0)(4)(47) xor ((not pi_in(1)(0)(47)) and pi_in(2)(1)(47));
 chi_out(3)(0)(48) <= pi_in(0)(4)(48) xor ((not pi_in(1)(0)(48)) and pi_in(2)(1)(48));
 chi_out(3)(0)(49) <= pi_in(0)(4)(49) xor ((not pi_in(1)(0)(49)) and pi_in(2)(1)(49));
 chi_out(3)(0)(50) <= pi_in(0)(4)(50) xor ((not pi_in(1)(0)(50)) and pi_in(2)(1)(50));
 chi_out(3)(0)(51) <= pi_in(0)(4)(51) xor ((not pi_in(1)(0)(51)) and pi_in(2)(1)(51));
 chi_out(3)(0)(52) <= pi_in(0)(4)(52) xor ((not pi_in(1)(0)(52)) and pi_in(2)(1)(52));
 chi_out(3)(0)(53) <= pi_in(0)(4)(53) xor ((not pi_in(1)(0)(53)) and pi_in(2)(1)(53));
 chi_out(3)(0)(54) <= pi_in(0)(4)(54) xor ((not pi_in(1)(0)(54)) and pi_in(2)(1)(54));
 chi_out(3)(0)(55) <= pi_in(0)(4)(55) xor ((not pi_in(1)(0)(55)) and pi_in(2)(1)(55));
 chi_out(3)(0)(56) <= pi_in(0)(4)(56) xor ((not pi_in(1)(0)(56)) and pi_in(2)(1)(56));
 chi_out(3)(0)(57) <= pi_in(0)(4)(57) xor ((not pi_in(1)(0)(57)) and pi_in(2)(1)(57));
 chi_out(3)(0)(58) <= pi_in(0)(4)(58) xor ((not pi_in(1)(0)(58)) and pi_in(2)(1)(58));
 chi_out(3)(0)(59) <= pi_in(0)(4)(59) xor ((not pi_in(1)(0)(59)) and pi_in(2)(1)(59));
 chi_out(3)(0)(60) <= pi_in(0)(4)(60) xor ((not pi_in(1)(0)(60)) and pi_in(2)(1)(60));
 chi_out(3)(0)(61) <= pi_in(0)(4)(61) xor ((not pi_in(1)(0)(61)) and pi_in(2)(1)(61));
 chi_out(3)(0)(62) <= pi_in(0)(4)(62) xor ((not pi_in(1)(0)(62)) and pi_in(2)(1)(62));
 chi_out(3)(0)(63) <= pi_in(0)(4)(63) xor ((not pi_in(1)(0)(63)) and pi_in(2)(1)(63));
 chi_out(3)(1)(0) <= pi_in(1)(0)(0) xor ((not pi_in(2)(1)(0)) and pi_in(3)(2)(0));
 chi_out(3)(1)(1) <= pi_in(1)(0)(1) xor ((not pi_in(2)(1)(1)) and pi_in(3)(2)(1));
 chi_out(3)(1)(2) <= pi_in(1)(0)(2) xor ((not pi_in(2)(1)(2)) and pi_in(3)(2)(2));
 chi_out(3)(1)(3) <= pi_in(1)(0)(3) xor ((not pi_in(2)(1)(3)) and pi_in(3)(2)(3));
 chi_out(3)(1)(4) <= pi_in(1)(0)(4) xor ((not pi_in(2)(1)(4)) and pi_in(3)(2)(4));
 chi_out(3)(1)(5) <= pi_in(1)(0)(5) xor ((not pi_in(2)(1)(5)) and pi_in(3)(2)(5));
 chi_out(3)(1)(6) <= pi_in(1)(0)(6) xor ((not pi_in(2)(1)(6)) and pi_in(3)(2)(6));
 chi_out(3)(1)(7) <= pi_in(1)(0)(7) xor ((not pi_in(2)(1)(7)) and pi_in(3)(2)(7));
 chi_out(3)(1)(8) <= pi_in(1)(0)(8) xor ((not pi_in(2)(1)(8)) and pi_in(3)(2)(8));
 chi_out(3)(1)(9) <= pi_in(1)(0)(9) xor ((not pi_in(2)(1)(9)) and pi_in(3)(2)(9));
 chi_out(3)(1)(10) <= pi_in(1)(0)(10) xor ((not pi_in(2)(1)(10)) and pi_in(3)(2)(10));
 chi_out(3)(1)(11) <= pi_in(1)(0)(11) xor ((not pi_in(2)(1)(11)) and pi_in(3)(2)(11));
 chi_out(3)(1)(12) <= pi_in(1)(0)(12) xor ((not pi_in(2)(1)(12)) and pi_in(3)(2)(12));
 chi_out(3)(1)(13) <= pi_in(1)(0)(13) xor ((not pi_in(2)(1)(13)) and pi_in(3)(2)(13));
 chi_out(3)(1)(14) <= pi_in(1)(0)(14) xor ((not pi_in(2)(1)(14)) and pi_in(3)(2)(14));
 chi_out(3)(1)(15) <= pi_in(1)(0)(15) xor ((not pi_in(2)(1)(15)) and pi_in(3)(2)(15));
 chi_out(3)(1)(16) <= pi_in(1)(0)(16) xor ((not pi_in(2)(1)(16)) and pi_in(3)(2)(16));
 chi_out(3)(1)(17) <= pi_in(1)(0)(17) xor ((not pi_in(2)(1)(17)) and pi_in(3)(2)(17));
 chi_out(3)(1)(18) <= pi_in(1)(0)(18) xor ((not pi_in(2)(1)(18)) and pi_in(3)(2)(18));
 chi_out(3)(1)(19) <= pi_in(1)(0)(19) xor ((not pi_in(2)(1)(19)) and pi_in(3)(2)(19));
 chi_out(3)(1)(20) <= pi_in(1)(0)(20) xor ((not pi_in(2)(1)(20)) and pi_in(3)(2)(20));
 chi_out(3)(1)(21) <= pi_in(1)(0)(21) xor ((not pi_in(2)(1)(21)) and pi_in(3)(2)(21));
 chi_out(3)(1)(22) <= pi_in(1)(0)(22) xor ((not pi_in(2)(1)(22)) and pi_in(3)(2)(22));
 chi_out(3)(1)(23) <= pi_in(1)(0)(23) xor ((not pi_in(2)(1)(23)) and pi_in(3)(2)(23));
 chi_out(3)(1)(24) <= pi_in(1)(0)(24) xor ((not pi_in(2)(1)(24)) and pi_in(3)(2)(24));
 chi_out(3)(1)(25) <= pi_in(1)(0)(25) xor ((not pi_in(2)(1)(25)) and pi_in(3)(2)(25));
 chi_out(3)(1)(26) <= pi_in(1)(0)(26) xor ((not pi_in(2)(1)(26)) and pi_in(3)(2)(26));
 chi_out(3)(1)(27) <= pi_in(1)(0)(27) xor ((not pi_in(2)(1)(27)) and pi_in(3)(2)(27));
 chi_out(3)(1)(28) <= pi_in(1)(0)(28) xor ((not pi_in(2)(1)(28)) and pi_in(3)(2)(28));
 chi_out(3)(1)(29) <= pi_in(1)(0)(29) xor ((not pi_in(2)(1)(29)) and pi_in(3)(2)(29));
 chi_out(3)(1)(30) <= pi_in(1)(0)(30) xor ((not pi_in(2)(1)(30)) and pi_in(3)(2)(30));
 chi_out(3)(1)(31) <= pi_in(1)(0)(31) xor ((not pi_in(2)(1)(31)) and pi_in(3)(2)(31));
 chi_out(3)(1)(32) <= pi_in(1)(0)(32) xor ((not pi_in(2)(1)(32)) and pi_in(3)(2)(32));
 chi_out(3)(1)(33) <= pi_in(1)(0)(33) xor ((not pi_in(2)(1)(33)) and pi_in(3)(2)(33));
 chi_out(3)(1)(34) <= pi_in(1)(0)(34) xor ((not pi_in(2)(1)(34)) and pi_in(3)(2)(34));
 chi_out(3)(1)(35) <= pi_in(1)(0)(35) xor ((not pi_in(2)(1)(35)) and pi_in(3)(2)(35));
 chi_out(3)(1)(36) <= pi_in(1)(0)(36) xor ((not pi_in(2)(1)(36)) and pi_in(3)(2)(36));
 chi_out(3)(1)(37) <= pi_in(1)(0)(37) xor ((not pi_in(2)(1)(37)) and pi_in(3)(2)(37));
 chi_out(3)(1)(38) <= pi_in(1)(0)(38) xor ((not pi_in(2)(1)(38)) and pi_in(3)(2)(38));
 chi_out(3)(1)(39) <= pi_in(1)(0)(39) xor ((not pi_in(2)(1)(39)) and pi_in(3)(2)(39));
 chi_out(3)(1)(40) <= pi_in(1)(0)(40) xor ((not pi_in(2)(1)(40)) and pi_in(3)(2)(40));
 chi_out(3)(1)(41) <= pi_in(1)(0)(41) xor ((not pi_in(2)(1)(41)) and pi_in(3)(2)(41));
 chi_out(3)(1)(42) <= pi_in(1)(0)(42) xor ((not pi_in(2)(1)(42)) and pi_in(3)(2)(42));
 chi_out(3)(1)(43) <= pi_in(1)(0)(43) xor ((not pi_in(2)(1)(43)) and pi_in(3)(2)(43));
 chi_out(3)(1)(44) <= pi_in(1)(0)(44) xor ((not pi_in(2)(1)(44)) and pi_in(3)(2)(44));
 chi_out(3)(1)(45) <= pi_in(1)(0)(45) xor ((not pi_in(2)(1)(45)) and pi_in(3)(2)(45));
 chi_out(3)(1)(46) <= pi_in(1)(0)(46) xor ((not pi_in(2)(1)(46)) and pi_in(3)(2)(46));
 chi_out(3)(1)(47) <= pi_in(1)(0)(47) xor ((not pi_in(2)(1)(47)) and pi_in(3)(2)(47));
 chi_out(3)(1)(48) <= pi_in(1)(0)(48) xor ((not pi_in(2)(1)(48)) and pi_in(3)(2)(48));
 chi_out(3)(1)(49) <= pi_in(1)(0)(49) xor ((not pi_in(2)(1)(49)) and pi_in(3)(2)(49));
 chi_out(3)(1)(50) <= pi_in(1)(0)(50) xor ((not pi_in(2)(1)(50)) and pi_in(3)(2)(50));
 chi_out(3)(1)(51) <= pi_in(1)(0)(51) xor ((not pi_in(2)(1)(51)) and pi_in(3)(2)(51));
 chi_out(3)(1)(52) <= pi_in(1)(0)(52) xor ((not pi_in(2)(1)(52)) and pi_in(3)(2)(52));
 chi_out(3)(1)(53) <= pi_in(1)(0)(53) xor ((not pi_in(2)(1)(53)) and pi_in(3)(2)(53));
 chi_out(3)(1)(54) <= pi_in(1)(0)(54) xor ((not pi_in(2)(1)(54)) and pi_in(3)(2)(54));
 chi_out(3)(1)(55) <= pi_in(1)(0)(55) xor ((not pi_in(2)(1)(55)) and pi_in(3)(2)(55));
 chi_out(3)(1)(56) <= pi_in(1)(0)(56) xor ((not pi_in(2)(1)(56)) and pi_in(3)(2)(56));
 chi_out(3)(1)(57) <= pi_in(1)(0)(57) xor ((not pi_in(2)(1)(57)) and pi_in(3)(2)(57));
 chi_out(3)(1)(58) <= pi_in(1)(0)(58) xor ((not pi_in(2)(1)(58)) and pi_in(3)(2)(58));
 chi_out(3)(1)(59) <= pi_in(1)(0)(59) xor ((not pi_in(2)(1)(59)) and pi_in(3)(2)(59));
 chi_out(3)(1)(60) <= pi_in(1)(0)(60) xor ((not pi_in(2)(1)(60)) and pi_in(3)(2)(60));
 chi_out(3)(1)(61) <= pi_in(1)(0)(61) xor ((not pi_in(2)(1)(61)) and pi_in(3)(2)(61));
 chi_out(3)(1)(62) <= pi_in(1)(0)(62) xor ((not pi_in(2)(1)(62)) and pi_in(3)(2)(62));
 chi_out(3)(1)(63) <= pi_in(1)(0)(63) xor ((not pi_in(2)(1)(63)) and pi_in(3)(2)(63));
 chi_out(3)(2)(0) <= pi_in(2)(1)(0) xor ((not pi_in(3)(2)(0)) and pi_in(4)(3)(0));
 chi_out(3)(2)(1) <= pi_in(2)(1)(1) xor ((not pi_in(3)(2)(1)) and pi_in(4)(3)(1));
 chi_out(3)(2)(2) <= pi_in(2)(1)(2) xor ((not pi_in(3)(2)(2)) and pi_in(4)(3)(2));
 chi_out(3)(2)(3) <= pi_in(2)(1)(3) xor ((not pi_in(3)(2)(3)) and pi_in(4)(3)(3));
 chi_out(3)(2)(4) <= pi_in(2)(1)(4) xor ((not pi_in(3)(2)(4)) and pi_in(4)(3)(4));
 chi_out(3)(2)(5) <= pi_in(2)(1)(5) xor ((not pi_in(3)(2)(5)) and pi_in(4)(3)(5));
 chi_out(3)(2)(6) <= pi_in(2)(1)(6) xor ((not pi_in(3)(2)(6)) and pi_in(4)(3)(6));
 chi_out(3)(2)(7) <= pi_in(2)(1)(7) xor ((not pi_in(3)(2)(7)) and pi_in(4)(3)(7));
 chi_out(3)(2)(8) <= pi_in(2)(1)(8) xor ((not pi_in(3)(2)(8)) and pi_in(4)(3)(8));
 chi_out(3)(2)(9) <= pi_in(2)(1)(9) xor ((not pi_in(3)(2)(9)) and pi_in(4)(3)(9));
 chi_out(3)(2)(10) <= pi_in(2)(1)(10) xor ((not pi_in(3)(2)(10)) and pi_in(4)(3)(10));
 chi_out(3)(2)(11) <= pi_in(2)(1)(11) xor ((not pi_in(3)(2)(11)) and pi_in(4)(3)(11));
 chi_out(3)(2)(12) <= pi_in(2)(1)(12) xor ((not pi_in(3)(2)(12)) and pi_in(4)(3)(12));
 chi_out(3)(2)(13) <= pi_in(2)(1)(13) xor ((not pi_in(3)(2)(13)) and pi_in(4)(3)(13));
 chi_out(3)(2)(14) <= pi_in(2)(1)(14) xor ((not pi_in(3)(2)(14)) and pi_in(4)(3)(14));
 chi_out(3)(2)(15) <= pi_in(2)(1)(15) xor ((not pi_in(3)(2)(15)) and pi_in(4)(3)(15));
 chi_out(3)(2)(16) <= pi_in(2)(1)(16) xor ((not pi_in(3)(2)(16)) and pi_in(4)(3)(16));
 chi_out(3)(2)(17) <= pi_in(2)(1)(17) xor ((not pi_in(3)(2)(17)) and pi_in(4)(3)(17));
 chi_out(3)(2)(18) <= pi_in(2)(1)(18) xor ((not pi_in(3)(2)(18)) and pi_in(4)(3)(18));
 chi_out(3)(2)(19) <= pi_in(2)(1)(19) xor ((not pi_in(3)(2)(19)) and pi_in(4)(3)(19));
 chi_out(3)(2)(20) <= pi_in(2)(1)(20) xor ((not pi_in(3)(2)(20)) and pi_in(4)(3)(20));
 chi_out(3)(2)(21) <= pi_in(2)(1)(21) xor ((not pi_in(3)(2)(21)) and pi_in(4)(3)(21));
 chi_out(3)(2)(22) <= pi_in(2)(1)(22) xor ((not pi_in(3)(2)(22)) and pi_in(4)(3)(22));
 chi_out(3)(2)(23) <= pi_in(2)(1)(23) xor ((not pi_in(3)(2)(23)) and pi_in(4)(3)(23));
 chi_out(3)(2)(24) <= pi_in(2)(1)(24) xor ((not pi_in(3)(2)(24)) and pi_in(4)(3)(24));
 chi_out(3)(2)(25) <= pi_in(2)(1)(25) xor ((not pi_in(3)(2)(25)) and pi_in(4)(3)(25));
 chi_out(3)(2)(26) <= pi_in(2)(1)(26) xor ((not pi_in(3)(2)(26)) and pi_in(4)(3)(26));
 chi_out(3)(2)(27) <= pi_in(2)(1)(27) xor ((not pi_in(3)(2)(27)) and pi_in(4)(3)(27));
 chi_out(3)(2)(28) <= pi_in(2)(1)(28) xor ((not pi_in(3)(2)(28)) and pi_in(4)(3)(28));
 chi_out(3)(2)(29) <= pi_in(2)(1)(29) xor ((not pi_in(3)(2)(29)) and pi_in(4)(3)(29));
 chi_out(3)(2)(30) <= pi_in(2)(1)(30) xor ((not pi_in(3)(2)(30)) and pi_in(4)(3)(30));
 chi_out(3)(2)(31) <= pi_in(2)(1)(31) xor ((not pi_in(3)(2)(31)) and pi_in(4)(3)(31));
 chi_out(3)(2)(32) <= pi_in(2)(1)(32) xor ((not pi_in(3)(2)(32)) and pi_in(4)(3)(32));
 chi_out(3)(2)(33) <= pi_in(2)(1)(33) xor ((not pi_in(3)(2)(33)) and pi_in(4)(3)(33));
 chi_out(3)(2)(34) <= pi_in(2)(1)(34) xor ((not pi_in(3)(2)(34)) and pi_in(4)(3)(34));
 chi_out(3)(2)(35) <= pi_in(2)(1)(35) xor ((not pi_in(3)(2)(35)) and pi_in(4)(3)(35));
 chi_out(3)(2)(36) <= pi_in(2)(1)(36) xor ((not pi_in(3)(2)(36)) and pi_in(4)(3)(36));
 chi_out(3)(2)(37) <= pi_in(2)(1)(37) xor ((not pi_in(3)(2)(37)) and pi_in(4)(3)(37));
 chi_out(3)(2)(38) <= pi_in(2)(1)(38) xor ((not pi_in(3)(2)(38)) and pi_in(4)(3)(38));
 chi_out(3)(2)(39) <= pi_in(2)(1)(39) xor ((not pi_in(3)(2)(39)) and pi_in(4)(3)(39));
 chi_out(3)(2)(40) <= pi_in(2)(1)(40) xor ((not pi_in(3)(2)(40)) and pi_in(4)(3)(40));
 chi_out(3)(2)(41) <= pi_in(2)(1)(41) xor ((not pi_in(3)(2)(41)) and pi_in(4)(3)(41));
 chi_out(3)(2)(42) <= pi_in(2)(1)(42) xor ((not pi_in(3)(2)(42)) and pi_in(4)(3)(42));
 chi_out(3)(2)(43) <= pi_in(2)(1)(43) xor ((not pi_in(3)(2)(43)) and pi_in(4)(3)(43));
 chi_out(3)(2)(44) <= pi_in(2)(1)(44) xor ((not pi_in(3)(2)(44)) and pi_in(4)(3)(44));
 chi_out(3)(2)(45) <= pi_in(2)(1)(45) xor ((not pi_in(3)(2)(45)) and pi_in(4)(3)(45));
 chi_out(3)(2)(46) <= pi_in(2)(1)(46) xor ((not pi_in(3)(2)(46)) and pi_in(4)(3)(46));
 chi_out(3)(2)(47) <= pi_in(2)(1)(47) xor ((not pi_in(3)(2)(47)) and pi_in(4)(3)(47));
 chi_out(3)(2)(48) <= pi_in(2)(1)(48) xor ((not pi_in(3)(2)(48)) and pi_in(4)(3)(48));
 chi_out(3)(2)(49) <= pi_in(2)(1)(49) xor ((not pi_in(3)(2)(49)) and pi_in(4)(3)(49));
 chi_out(3)(2)(50) <= pi_in(2)(1)(50) xor ((not pi_in(3)(2)(50)) and pi_in(4)(3)(50));
 chi_out(3)(2)(51) <= pi_in(2)(1)(51) xor ((not pi_in(3)(2)(51)) and pi_in(4)(3)(51));
 chi_out(3)(2)(52) <= pi_in(2)(1)(52) xor ((not pi_in(3)(2)(52)) and pi_in(4)(3)(52));
 chi_out(3)(2)(53) <= pi_in(2)(1)(53) xor ((not pi_in(3)(2)(53)) and pi_in(4)(3)(53));
 chi_out(3)(2)(54) <= pi_in(2)(1)(54) xor ((not pi_in(3)(2)(54)) and pi_in(4)(3)(54));
 chi_out(3)(2)(55) <= pi_in(2)(1)(55) xor ((not pi_in(3)(2)(55)) and pi_in(4)(3)(55));
 chi_out(3)(2)(56) <= pi_in(2)(1)(56) xor ((not pi_in(3)(2)(56)) and pi_in(4)(3)(56));
 chi_out(3)(2)(57) <= pi_in(2)(1)(57) xor ((not pi_in(3)(2)(57)) and pi_in(4)(3)(57));
 chi_out(3)(2)(58) <= pi_in(2)(1)(58) xor ((not pi_in(3)(2)(58)) and pi_in(4)(3)(58));
 chi_out(3)(2)(59) <= pi_in(2)(1)(59) xor ((not pi_in(3)(2)(59)) and pi_in(4)(3)(59));
 chi_out(3)(2)(60) <= pi_in(2)(1)(60) xor ((not pi_in(3)(2)(60)) and pi_in(4)(3)(60));
 chi_out(3)(2)(61) <= pi_in(2)(1)(61) xor ((not pi_in(3)(2)(61)) and pi_in(4)(3)(61));
 chi_out(3)(2)(62) <= pi_in(2)(1)(62) xor ((not pi_in(3)(2)(62)) and pi_in(4)(3)(62));
 chi_out(3)(2)(63) <= pi_in(2)(1)(63) xor ((not pi_in(3)(2)(63)) and pi_in(4)(3)(63));
 chi_out(4)(0)(0) <= pi_in(0)(2)(0) xor ((not pi_in(1)(3)(0)) and pi_in(2)(4)(0));
 chi_out(4)(0)(1) <= pi_in(0)(2)(1) xor ((not pi_in(1)(3)(1)) and pi_in(2)(4)(1));
 chi_out(4)(0)(2) <= pi_in(0)(2)(2) xor ((not pi_in(1)(3)(2)) and pi_in(2)(4)(2));
 chi_out(4)(0)(3) <= pi_in(0)(2)(3) xor ((not pi_in(1)(3)(3)) and pi_in(2)(4)(3));
 chi_out(4)(0)(4) <= pi_in(0)(2)(4) xor ((not pi_in(1)(3)(4)) and pi_in(2)(4)(4));
 chi_out(4)(0)(5) <= pi_in(0)(2)(5) xor ((not pi_in(1)(3)(5)) and pi_in(2)(4)(5));
 chi_out(4)(0)(6) <= pi_in(0)(2)(6) xor ((not pi_in(1)(3)(6)) and pi_in(2)(4)(6));
 chi_out(4)(0)(7) <= pi_in(0)(2)(7) xor ((not pi_in(1)(3)(7)) and pi_in(2)(4)(7));
 chi_out(4)(0)(8) <= pi_in(0)(2)(8) xor ((not pi_in(1)(3)(8)) and pi_in(2)(4)(8));
 chi_out(4)(0)(9) <= pi_in(0)(2)(9) xor ((not pi_in(1)(3)(9)) and pi_in(2)(4)(9));
 chi_out(4)(0)(10) <= pi_in(0)(2)(10) xor ((not pi_in(1)(3)(10)) and pi_in(2)(4)(10));
 chi_out(4)(0)(11) <= pi_in(0)(2)(11) xor ((not pi_in(1)(3)(11)) and pi_in(2)(4)(11));
 chi_out(4)(0)(12) <= pi_in(0)(2)(12) xor ((not pi_in(1)(3)(12)) and pi_in(2)(4)(12));
 chi_out(4)(0)(13) <= pi_in(0)(2)(13) xor ((not pi_in(1)(3)(13)) and pi_in(2)(4)(13));
 chi_out(4)(0)(14) <= pi_in(0)(2)(14) xor ((not pi_in(1)(3)(14)) and pi_in(2)(4)(14));
 chi_out(4)(0)(15) <= pi_in(0)(2)(15) xor ((not pi_in(1)(3)(15)) and pi_in(2)(4)(15));
 chi_out(4)(0)(16) <= pi_in(0)(2)(16) xor ((not pi_in(1)(3)(16)) and pi_in(2)(4)(16));
 chi_out(4)(0)(17) <= pi_in(0)(2)(17) xor ((not pi_in(1)(3)(17)) and pi_in(2)(4)(17));
 chi_out(4)(0)(18) <= pi_in(0)(2)(18) xor ((not pi_in(1)(3)(18)) and pi_in(2)(4)(18));
 chi_out(4)(0)(19) <= pi_in(0)(2)(19) xor ((not pi_in(1)(3)(19)) and pi_in(2)(4)(19));
 chi_out(4)(0)(20) <= pi_in(0)(2)(20) xor ((not pi_in(1)(3)(20)) and pi_in(2)(4)(20));
 chi_out(4)(0)(21) <= pi_in(0)(2)(21) xor ((not pi_in(1)(3)(21)) and pi_in(2)(4)(21));
 chi_out(4)(0)(22) <= pi_in(0)(2)(22) xor ((not pi_in(1)(3)(22)) and pi_in(2)(4)(22));
 chi_out(4)(0)(23) <= pi_in(0)(2)(23) xor ((not pi_in(1)(3)(23)) and pi_in(2)(4)(23));
 chi_out(4)(0)(24) <= pi_in(0)(2)(24) xor ((not pi_in(1)(3)(24)) and pi_in(2)(4)(24));
 chi_out(4)(0)(25) <= pi_in(0)(2)(25) xor ((not pi_in(1)(3)(25)) and pi_in(2)(4)(25));
 chi_out(4)(0)(26) <= pi_in(0)(2)(26) xor ((not pi_in(1)(3)(26)) and pi_in(2)(4)(26));
 chi_out(4)(0)(27) <= pi_in(0)(2)(27) xor ((not pi_in(1)(3)(27)) and pi_in(2)(4)(27));
 chi_out(4)(0)(28) <= pi_in(0)(2)(28) xor ((not pi_in(1)(3)(28)) and pi_in(2)(4)(28));
 chi_out(4)(0)(29) <= pi_in(0)(2)(29) xor ((not pi_in(1)(3)(29)) and pi_in(2)(4)(29));
 chi_out(4)(0)(30) <= pi_in(0)(2)(30) xor ((not pi_in(1)(3)(30)) and pi_in(2)(4)(30));
 chi_out(4)(0)(31) <= pi_in(0)(2)(31) xor ((not pi_in(1)(3)(31)) and pi_in(2)(4)(31));
 chi_out(4)(0)(32) <= pi_in(0)(2)(32) xor ((not pi_in(1)(3)(32)) and pi_in(2)(4)(32));
 chi_out(4)(0)(33) <= pi_in(0)(2)(33) xor ((not pi_in(1)(3)(33)) and pi_in(2)(4)(33));
 chi_out(4)(0)(34) <= pi_in(0)(2)(34) xor ((not pi_in(1)(3)(34)) and pi_in(2)(4)(34));
 chi_out(4)(0)(35) <= pi_in(0)(2)(35) xor ((not pi_in(1)(3)(35)) and pi_in(2)(4)(35));
 chi_out(4)(0)(36) <= pi_in(0)(2)(36) xor ((not pi_in(1)(3)(36)) and pi_in(2)(4)(36));
 chi_out(4)(0)(37) <= pi_in(0)(2)(37) xor ((not pi_in(1)(3)(37)) and pi_in(2)(4)(37));
 chi_out(4)(0)(38) <= pi_in(0)(2)(38) xor ((not pi_in(1)(3)(38)) and pi_in(2)(4)(38));
 chi_out(4)(0)(39) <= pi_in(0)(2)(39) xor ((not pi_in(1)(3)(39)) and pi_in(2)(4)(39));
 chi_out(4)(0)(40) <= pi_in(0)(2)(40) xor ((not pi_in(1)(3)(40)) and pi_in(2)(4)(40));
 chi_out(4)(0)(41) <= pi_in(0)(2)(41) xor ((not pi_in(1)(3)(41)) and pi_in(2)(4)(41));
 chi_out(4)(0)(42) <= pi_in(0)(2)(42) xor ((not pi_in(1)(3)(42)) and pi_in(2)(4)(42));
 chi_out(4)(0)(43) <= pi_in(0)(2)(43) xor ((not pi_in(1)(3)(43)) and pi_in(2)(4)(43));
 chi_out(4)(0)(44) <= pi_in(0)(2)(44) xor ((not pi_in(1)(3)(44)) and pi_in(2)(4)(44));
 chi_out(4)(0)(45) <= pi_in(0)(2)(45) xor ((not pi_in(1)(3)(45)) and pi_in(2)(4)(45));
 chi_out(4)(0)(46) <= pi_in(0)(2)(46) xor ((not pi_in(1)(3)(46)) and pi_in(2)(4)(46));
 chi_out(4)(0)(47) <= pi_in(0)(2)(47) xor ((not pi_in(1)(3)(47)) and pi_in(2)(4)(47));
 chi_out(4)(0)(48) <= pi_in(0)(2)(48) xor ((not pi_in(1)(3)(48)) and pi_in(2)(4)(48));
 chi_out(4)(0)(49) <= pi_in(0)(2)(49) xor ((not pi_in(1)(3)(49)) and pi_in(2)(4)(49));
 chi_out(4)(0)(50) <= pi_in(0)(2)(50) xor ((not pi_in(1)(3)(50)) and pi_in(2)(4)(50));
 chi_out(4)(0)(51) <= pi_in(0)(2)(51) xor ((not pi_in(1)(3)(51)) and pi_in(2)(4)(51));
 chi_out(4)(0)(52) <= pi_in(0)(2)(52) xor ((not pi_in(1)(3)(52)) and pi_in(2)(4)(52));
 chi_out(4)(0)(53) <= pi_in(0)(2)(53) xor ((not pi_in(1)(3)(53)) and pi_in(2)(4)(53));
 chi_out(4)(0)(54) <= pi_in(0)(2)(54) xor ((not pi_in(1)(3)(54)) and pi_in(2)(4)(54));
 chi_out(4)(0)(55) <= pi_in(0)(2)(55) xor ((not pi_in(1)(3)(55)) and pi_in(2)(4)(55));
 chi_out(4)(0)(56) <= pi_in(0)(2)(56) xor ((not pi_in(1)(3)(56)) and pi_in(2)(4)(56));
 chi_out(4)(0)(57) <= pi_in(0)(2)(57) xor ((not pi_in(1)(3)(57)) and pi_in(2)(4)(57));
 chi_out(4)(0)(58) <= pi_in(0)(2)(58) xor ((not pi_in(1)(3)(58)) and pi_in(2)(4)(58));
 chi_out(4)(0)(59) <= pi_in(0)(2)(59) xor ((not pi_in(1)(3)(59)) and pi_in(2)(4)(59));
 chi_out(4)(0)(60) <= pi_in(0)(2)(60) xor ((not pi_in(1)(3)(60)) and pi_in(2)(4)(60));
 chi_out(4)(0)(61) <= pi_in(0)(2)(61) xor ((not pi_in(1)(3)(61)) and pi_in(2)(4)(61));
 chi_out(4)(0)(62) <= pi_in(0)(2)(62) xor ((not pi_in(1)(3)(62)) and pi_in(2)(4)(62));
 chi_out(4)(0)(63) <= pi_in(0)(2)(63) xor ((not pi_in(1)(3)(63)) and pi_in(2)(4)(63));
 chi_out(4)(1)(0) <= pi_in(1)(3)(0) xor ((not pi_in(2)(4)(0)) and pi_in(3)(0)(0));
 chi_out(4)(1)(1) <= pi_in(1)(3)(1) xor ((not pi_in(2)(4)(1)) and pi_in(3)(0)(1));
 chi_out(4)(1)(2) <= pi_in(1)(3)(2) xor ((not pi_in(2)(4)(2)) and pi_in(3)(0)(2));
 chi_out(4)(1)(3) <= pi_in(1)(3)(3) xor ((not pi_in(2)(4)(3)) and pi_in(3)(0)(3));
 chi_out(4)(1)(4) <= pi_in(1)(3)(4) xor ((not pi_in(2)(4)(4)) and pi_in(3)(0)(4));
 chi_out(4)(1)(5) <= pi_in(1)(3)(5) xor ((not pi_in(2)(4)(5)) and pi_in(3)(0)(5));
 chi_out(4)(1)(6) <= pi_in(1)(3)(6) xor ((not pi_in(2)(4)(6)) and pi_in(3)(0)(6));
 chi_out(4)(1)(7) <= pi_in(1)(3)(7) xor ((not pi_in(2)(4)(7)) and pi_in(3)(0)(7));
 chi_out(4)(1)(8) <= pi_in(1)(3)(8) xor ((not pi_in(2)(4)(8)) and pi_in(3)(0)(8));
 chi_out(4)(1)(9) <= pi_in(1)(3)(9) xor ((not pi_in(2)(4)(9)) and pi_in(3)(0)(9));
 chi_out(4)(1)(10) <= pi_in(1)(3)(10) xor ((not pi_in(2)(4)(10)) and pi_in(3)(0)(10));
 chi_out(4)(1)(11) <= pi_in(1)(3)(11) xor ((not pi_in(2)(4)(11)) and pi_in(3)(0)(11));
 chi_out(4)(1)(12) <= pi_in(1)(3)(12) xor ((not pi_in(2)(4)(12)) and pi_in(3)(0)(12));
 chi_out(4)(1)(13) <= pi_in(1)(3)(13) xor ((not pi_in(2)(4)(13)) and pi_in(3)(0)(13));
 chi_out(4)(1)(14) <= pi_in(1)(3)(14) xor ((not pi_in(2)(4)(14)) and pi_in(3)(0)(14));
 chi_out(4)(1)(15) <= pi_in(1)(3)(15) xor ((not pi_in(2)(4)(15)) and pi_in(3)(0)(15));
 chi_out(4)(1)(16) <= pi_in(1)(3)(16) xor ((not pi_in(2)(4)(16)) and pi_in(3)(0)(16));
 chi_out(4)(1)(17) <= pi_in(1)(3)(17) xor ((not pi_in(2)(4)(17)) and pi_in(3)(0)(17));
 chi_out(4)(1)(18) <= pi_in(1)(3)(18) xor ((not pi_in(2)(4)(18)) and pi_in(3)(0)(18));
 chi_out(4)(1)(19) <= pi_in(1)(3)(19) xor ((not pi_in(2)(4)(19)) and pi_in(3)(0)(19));
 chi_out(4)(1)(20) <= pi_in(1)(3)(20) xor ((not pi_in(2)(4)(20)) and pi_in(3)(0)(20));
 chi_out(4)(1)(21) <= pi_in(1)(3)(21) xor ((not pi_in(2)(4)(21)) and pi_in(3)(0)(21));
 chi_out(4)(1)(22) <= pi_in(1)(3)(22) xor ((not pi_in(2)(4)(22)) and pi_in(3)(0)(22));
 chi_out(4)(1)(23) <= pi_in(1)(3)(23) xor ((not pi_in(2)(4)(23)) and pi_in(3)(0)(23));
 chi_out(4)(1)(24) <= pi_in(1)(3)(24) xor ((not pi_in(2)(4)(24)) and pi_in(3)(0)(24));
 chi_out(4)(1)(25) <= pi_in(1)(3)(25) xor ((not pi_in(2)(4)(25)) and pi_in(3)(0)(25));
 chi_out(4)(1)(26) <= pi_in(1)(3)(26) xor ((not pi_in(2)(4)(26)) and pi_in(3)(0)(26));
 chi_out(4)(1)(27) <= pi_in(1)(3)(27) xor ((not pi_in(2)(4)(27)) and pi_in(3)(0)(27));
 chi_out(4)(1)(28) <= pi_in(1)(3)(28) xor ((not pi_in(2)(4)(28)) and pi_in(3)(0)(28));
 chi_out(4)(1)(29) <= pi_in(1)(3)(29) xor ((not pi_in(2)(4)(29)) and pi_in(3)(0)(29));
 chi_out(4)(1)(30) <= pi_in(1)(3)(30) xor ((not pi_in(2)(4)(30)) and pi_in(3)(0)(30));
 chi_out(4)(1)(31) <= pi_in(1)(3)(31) xor ((not pi_in(2)(4)(31)) and pi_in(3)(0)(31));
 chi_out(4)(1)(32) <= pi_in(1)(3)(32) xor ((not pi_in(2)(4)(32)) and pi_in(3)(0)(32));
 chi_out(4)(1)(33) <= pi_in(1)(3)(33) xor ((not pi_in(2)(4)(33)) and pi_in(3)(0)(33));
 chi_out(4)(1)(34) <= pi_in(1)(3)(34) xor ((not pi_in(2)(4)(34)) and pi_in(3)(0)(34));
 chi_out(4)(1)(35) <= pi_in(1)(3)(35) xor ((not pi_in(2)(4)(35)) and pi_in(3)(0)(35));
 chi_out(4)(1)(36) <= pi_in(1)(3)(36) xor ((not pi_in(2)(4)(36)) and pi_in(3)(0)(36));
 chi_out(4)(1)(37) <= pi_in(1)(3)(37) xor ((not pi_in(2)(4)(37)) and pi_in(3)(0)(37));
 chi_out(4)(1)(38) <= pi_in(1)(3)(38) xor ((not pi_in(2)(4)(38)) and pi_in(3)(0)(38));
 chi_out(4)(1)(39) <= pi_in(1)(3)(39) xor ((not pi_in(2)(4)(39)) and pi_in(3)(0)(39));
 chi_out(4)(1)(40) <= pi_in(1)(3)(40) xor ((not pi_in(2)(4)(40)) and pi_in(3)(0)(40));
 chi_out(4)(1)(41) <= pi_in(1)(3)(41) xor ((not pi_in(2)(4)(41)) and pi_in(3)(0)(41));
 chi_out(4)(1)(42) <= pi_in(1)(3)(42) xor ((not pi_in(2)(4)(42)) and pi_in(3)(0)(42));
 chi_out(4)(1)(43) <= pi_in(1)(3)(43) xor ((not pi_in(2)(4)(43)) and pi_in(3)(0)(43));
 chi_out(4)(1)(44) <= pi_in(1)(3)(44) xor ((not pi_in(2)(4)(44)) and pi_in(3)(0)(44));
 chi_out(4)(1)(45) <= pi_in(1)(3)(45) xor ((not pi_in(2)(4)(45)) and pi_in(3)(0)(45));
 chi_out(4)(1)(46) <= pi_in(1)(3)(46) xor ((not pi_in(2)(4)(46)) and pi_in(3)(0)(46));
 chi_out(4)(1)(47) <= pi_in(1)(3)(47) xor ((not pi_in(2)(4)(47)) and pi_in(3)(0)(47));
 chi_out(4)(1)(48) <= pi_in(1)(3)(48) xor ((not pi_in(2)(4)(48)) and pi_in(3)(0)(48));
 chi_out(4)(1)(49) <= pi_in(1)(3)(49) xor ((not pi_in(2)(4)(49)) and pi_in(3)(0)(49));
 chi_out(4)(1)(50) <= pi_in(1)(3)(50) xor ((not pi_in(2)(4)(50)) and pi_in(3)(0)(50));
 chi_out(4)(1)(51) <= pi_in(1)(3)(51) xor ((not pi_in(2)(4)(51)) and pi_in(3)(0)(51));
 chi_out(4)(1)(52) <= pi_in(1)(3)(52) xor ((not pi_in(2)(4)(52)) and pi_in(3)(0)(52));
 chi_out(4)(1)(53) <= pi_in(1)(3)(53) xor ((not pi_in(2)(4)(53)) and pi_in(3)(0)(53));
 chi_out(4)(1)(54) <= pi_in(1)(3)(54) xor ((not pi_in(2)(4)(54)) and pi_in(3)(0)(54));
 chi_out(4)(1)(55) <= pi_in(1)(3)(55) xor ((not pi_in(2)(4)(55)) and pi_in(3)(0)(55));
 chi_out(4)(1)(56) <= pi_in(1)(3)(56) xor ((not pi_in(2)(4)(56)) and pi_in(3)(0)(56));
 chi_out(4)(1)(57) <= pi_in(1)(3)(57) xor ((not pi_in(2)(4)(57)) and pi_in(3)(0)(57));
 chi_out(4)(1)(58) <= pi_in(1)(3)(58) xor ((not pi_in(2)(4)(58)) and pi_in(3)(0)(58));
 chi_out(4)(1)(59) <= pi_in(1)(3)(59) xor ((not pi_in(2)(4)(59)) and pi_in(3)(0)(59));
 chi_out(4)(1)(60) <= pi_in(1)(3)(60) xor ((not pi_in(2)(4)(60)) and pi_in(3)(0)(60));
 chi_out(4)(1)(61) <= pi_in(1)(3)(61) xor ((not pi_in(2)(4)(61)) and pi_in(3)(0)(61));
 chi_out(4)(1)(62) <= pi_in(1)(3)(62) xor ((not pi_in(2)(4)(62)) and pi_in(3)(0)(62));
 chi_out(4)(1)(63) <= pi_in(1)(3)(63) xor ((not pi_in(2)(4)(63)) and pi_in(3)(0)(63));
 chi_out(4)(2)(0) <= pi_in(2)(4)(0) xor ((not pi_in(3)(0)(0)) and pi_in(4)(1)(0));
 chi_out(4)(2)(1) <= pi_in(2)(4)(1) xor ((not pi_in(3)(0)(1)) and pi_in(4)(1)(1));
 chi_out(4)(2)(2) <= pi_in(2)(4)(2) xor ((not pi_in(3)(0)(2)) and pi_in(4)(1)(2));
 chi_out(4)(2)(3) <= pi_in(2)(4)(3) xor ((not pi_in(3)(0)(3)) and pi_in(4)(1)(3));
 chi_out(4)(2)(4) <= pi_in(2)(4)(4) xor ((not pi_in(3)(0)(4)) and pi_in(4)(1)(4));
 chi_out(4)(2)(5) <= pi_in(2)(4)(5) xor ((not pi_in(3)(0)(5)) and pi_in(4)(1)(5));
 chi_out(4)(2)(6) <= pi_in(2)(4)(6) xor ((not pi_in(3)(0)(6)) and pi_in(4)(1)(6));
 chi_out(4)(2)(7) <= pi_in(2)(4)(7) xor ((not pi_in(3)(0)(7)) and pi_in(4)(1)(7));
 chi_out(4)(2)(8) <= pi_in(2)(4)(8) xor ((not pi_in(3)(0)(8)) and pi_in(4)(1)(8));
 chi_out(4)(2)(9) <= pi_in(2)(4)(9) xor ((not pi_in(3)(0)(9)) and pi_in(4)(1)(9));
 chi_out(4)(2)(10) <= pi_in(2)(4)(10) xor ((not pi_in(3)(0)(10)) and pi_in(4)(1)(10));
 chi_out(4)(2)(11) <= pi_in(2)(4)(11) xor ((not pi_in(3)(0)(11)) and pi_in(4)(1)(11));
 chi_out(4)(2)(12) <= pi_in(2)(4)(12) xor ((not pi_in(3)(0)(12)) and pi_in(4)(1)(12));
 chi_out(4)(2)(13) <= pi_in(2)(4)(13) xor ((not pi_in(3)(0)(13)) and pi_in(4)(1)(13));
 chi_out(4)(2)(14) <= pi_in(2)(4)(14) xor ((not pi_in(3)(0)(14)) and pi_in(4)(1)(14));
 chi_out(4)(2)(15) <= pi_in(2)(4)(15) xor ((not pi_in(3)(0)(15)) and pi_in(4)(1)(15));
 chi_out(4)(2)(16) <= pi_in(2)(4)(16) xor ((not pi_in(3)(0)(16)) and pi_in(4)(1)(16));
 chi_out(4)(2)(17) <= pi_in(2)(4)(17) xor ((not pi_in(3)(0)(17)) and pi_in(4)(1)(17));
 chi_out(4)(2)(18) <= pi_in(2)(4)(18) xor ((not pi_in(3)(0)(18)) and pi_in(4)(1)(18));
 chi_out(4)(2)(19) <= pi_in(2)(4)(19) xor ((not pi_in(3)(0)(19)) and pi_in(4)(1)(19));
 chi_out(4)(2)(20) <= pi_in(2)(4)(20) xor ((not pi_in(3)(0)(20)) and pi_in(4)(1)(20));
 chi_out(4)(2)(21) <= pi_in(2)(4)(21) xor ((not pi_in(3)(0)(21)) and pi_in(4)(1)(21));
 chi_out(4)(2)(22) <= pi_in(2)(4)(22) xor ((not pi_in(3)(0)(22)) and pi_in(4)(1)(22));
 chi_out(4)(2)(23) <= pi_in(2)(4)(23) xor ((not pi_in(3)(0)(23)) and pi_in(4)(1)(23));
 chi_out(4)(2)(24) <= pi_in(2)(4)(24) xor ((not pi_in(3)(0)(24)) and pi_in(4)(1)(24));
 chi_out(4)(2)(25) <= pi_in(2)(4)(25) xor ((not pi_in(3)(0)(25)) and pi_in(4)(1)(25));
 chi_out(4)(2)(26) <= pi_in(2)(4)(26) xor ((not pi_in(3)(0)(26)) and pi_in(4)(1)(26));
 chi_out(4)(2)(27) <= pi_in(2)(4)(27) xor ((not pi_in(3)(0)(27)) and pi_in(4)(1)(27));
 chi_out(4)(2)(28) <= pi_in(2)(4)(28) xor ((not pi_in(3)(0)(28)) and pi_in(4)(1)(28));
 chi_out(4)(2)(29) <= pi_in(2)(4)(29) xor ((not pi_in(3)(0)(29)) and pi_in(4)(1)(29));
 chi_out(4)(2)(30) <= pi_in(2)(4)(30) xor ((not pi_in(3)(0)(30)) and pi_in(4)(1)(30));
 chi_out(4)(2)(31) <= pi_in(2)(4)(31) xor ((not pi_in(3)(0)(31)) and pi_in(4)(1)(31));
 chi_out(4)(2)(32) <= pi_in(2)(4)(32) xor ((not pi_in(3)(0)(32)) and pi_in(4)(1)(32));
 chi_out(4)(2)(33) <= pi_in(2)(4)(33) xor ((not pi_in(3)(0)(33)) and pi_in(4)(1)(33));
 chi_out(4)(2)(34) <= pi_in(2)(4)(34) xor ((not pi_in(3)(0)(34)) and pi_in(4)(1)(34));
 chi_out(4)(2)(35) <= pi_in(2)(4)(35) xor ((not pi_in(3)(0)(35)) and pi_in(4)(1)(35));
 chi_out(4)(2)(36) <= pi_in(2)(4)(36) xor ((not pi_in(3)(0)(36)) and pi_in(4)(1)(36));
 chi_out(4)(2)(37) <= pi_in(2)(4)(37) xor ((not pi_in(3)(0)(37)) and pi_in(4)(1)(37));
 chi_out(4)(2)(38) <= pi_in(2)(4)(38) xor ((not pi_in(3)(0)(38)) and pi_in(4)(1)(38));
 chi_out(4)(2)(39) <= pi_in(2)(4)(39) xor ((not pi_in(3)(0)(39)) and pi_in(4)(1)(39));
 chi_out(4)(2)(40) <= pi_in(2)(4)(40) xor ((not pi_in(3)(0)(40)) and pi_in(4)(1)(40));
 chi_out(4)(2)(41) <= pi_in(2)(4)(41) xor ((not pi_in(3)(0)(41)) and pi_in(4)(1)(41));
 chi_out(4)(2)(42) <= pi_in(2)(4)(42) xor ((not pi_in(3)(0)(42)) and pi_in(4)(1)(42));
 chi_out(4)(2)(43) <= pi_in(2)(4)(43) xor ((not pi_in(3)(0)(43)) and pi_in(4)(1)(43));
 chi_out(4)(2)(44) <= pi_in(2)(4)(44) xor ((not pi_in(3)(0)(44)) and pi_in(4)(1)(44));
 chi_out(4)(2)(45) <= pi_in(2)(4)(45) xor ((not pi_in(3)(0)(45)) and pi_in(4)(1)(45));
 chi_out(4)(2)(46) <= pi_in(2)(4)(46) xor ((not pi_in(3)(0)(46)) and pi_in(4)(1)(46));
 chi_out(4)(2)(47) <= pi_in(2)(4)(47) xor ((not pi_in(3)(0)(47)) and pi_in(4)(1)(47));
 chi_out(4)(2)(48) <= pi_in(2)(4)(48) xor ((not pi_in(3)(0)(48)) and pi_in(4)(1)(48));
 chi_out(4)(2)(49) <= pi_in(2)(4)(49) xor ((not pi_in(3)(0)(49)) and pi_in(4)(1)(49));
 chi_out(4)(2)(50) <= pi_in(2)(4)(50) xor ((not pi_in(3)(0)(50)) and pi_in(4)(1)(50));
 chi_out(4)(2)(51) <= pi_in(2)(4)(51) xor ((not pi_in(3)(0)(51)) and pi_in(4)(1)(51));
 chi_out(4)(2)(52) <= pi_in(2)(4)(52) xor ((not pi_in(3)(0)(52)) and pi_in(4)(1)(52));
 chi_out(4)(2)(53) <= pi_in(2)(4)(53) xor ((not pi_in(3)(0)(53)) and pi_in(4)(1)(53));
 chi_out(4)(2)(54) <= pi_in(2)(4)(54) xor ((not pi_in(3)(0)(54)) and pi_in(4)(1)(54));
 chi_out(4)(2)(55) <= pi_in(2)(4)(55) xor ((not pi_in(3)(0)(55)) and pi_in(4)(1)(55));
 chi_out(4)(2)(56) <= pi_in(2)(4)(56) xor ((not pi_in(3)(0)(56)) and pi_in(4)(1)(56));
 chi_out(4)(2)(57) <= pi_in(2)(4)(57) xor ((not pi_in(3)(0)(57)) and pi_in(4)(1)(57));
 chi_out(4)(2)(58) <= pi_in(2)(4)(58) xor ((not pi_in(3)(0)(58)) and pi_in(4)(1)(58));
 chi_out(4)(2)(59) <= pi_in(2)(4)(59) xor ((not pi_in(3)(0)(59)) and pi_in(4)(1)(59));
 chi_out(4)(2)(60) <= pi_in(2)(4)(60) xor ((not pi_in(3)(0)(60)) and pi_in(4)(1)(60));
 chi_out(4)(2)(61) <= pi_in(2)(4)(61) xor ((not pi_in(3)(0)(61)) and pi_in(4)(1)(61));
 chi_out(4)(2)(62) <= pi_in(2)(4)(62) xor ((not pi_in(3)(0)(62)) and pi_in(4)(1)(62));
 chi_out(4)(2)(63) <= pi_in(2)(4)(63) xor ((not pi_in(3)(0)(63)) and pi_in(4)(1)(63));
 chi_out(0)(3)(0) <= pi_in(3)(3)(0) xor ((not pi_in(4)(4)(0)) and pi_in(0)(0)(0));
 chi_out(0)(3)(1) <= pi_in(3)(3)(1) xor ((not pi_in(4)(4)(1)) and pi_in(0)(0)(1));
 chi_out(0)(3)(2) <= pi_in(3)(3)(2) xor ((not pi_in(4)(4)(2)) and pi_in(0)(0)(2));
 chi_out(0)(3)(3) <= pi_in(3)(3)(3) xor ((not pi_in(4)(4)(3)) and pi_in(0)(0)(3));
 chi_out(0)(3)(4) <= pi_in(3)(3)(4) xor ((not pi_in(4)(4)(4)) and pi_in(0)(0)(4));
 chi_out(0)(3)(5) <= pi_in(3)(3)(5) xor ((not pi_in(4)(4)(5)) and pi_in(0)(0)(5));
 chi_out(0)(3)(6) <= pi_in(3)(3)(6) xor ((not pi_in(4)(4)(6)) and pi_in(0)(0)(6));
 chi_out(0)(3)(7) <= pi_in(3)(3)(7) xor ((not pi_in(4)(4)(7)) and pi_in(0)(0)(7));
 chi_out(0)(3)(8) <= pi_in(3)(3)(8) xor ((not pi_in(4)(4)(8)) and pi_in(0)(0)(8));
 chi_out(0)(3)(9) <= pi_in(3)(3)(9) xor ((not pi_in(4)(4)(9)) and pi_in(0)(0)(9));
 chi_out(0)(3)(10) <= pi_in(3)(3)(10) xor ((not pi_in(4)(4)(10)) and pi_in(0)(0)(10));
 chi_out(0)(3)(11) <= pi_in(3)(3)(11) xor ((not pi_in(4)(4)(11)) and pi_in(0)(0)(11));
 chi_out(0)(3)(12) <= pi_in(3)(3)(12) xor ((not pi_in(4)(4)(12)) and pi_in(0)(0)(12));
 chi_out(0)(3)(13) <= pi_in(3)(3)(13) xor ((not pi_in(4)(4)(13)) and pi_in(0)(0)(13));
 chi_out(0)(3)(14) <= pi_in(3)(3)(14) xor ((not pi_in(4)(4)(14)) and pi_in(0)(0)(14));
 chi_out(0)(3)(15) <= pi_in(3)(3)(15) xor ((not pi_in(4)(4)(15)) and pi_in(0)(0)(15));
 chi_out(0)(3)(16) <= pi_in(3)(3)(16) xor ((not pi_in(4)(4)(16)) and pi_in(0)(0)(16));
 chi_out(0)(3)(17) <= pi_in(3)(3)(17) xor ((not pi_in(4)(4)(17)) and pi_in(0)(0)(17));
 chi_out(0)(3)(18) <= pi_in(3)(3)(18) xor ((not pi_in(4)(4)(18)) and pi_in(0)(0)(18));
 chi_out(0)(3)(19) <= pi_in(3)(3)(19) xor ((not pi_in(4)(4)(19)) and pi_in(0)(0)(19));
 chi_out(0)(3)(20) <= pi_in(3)(3)(20) xor ((not pi_in(4)(4)(20)) and pi_in(0)(0)(20));
 chi_out(0)(3)(21) <= pi_in(3)(3)(21) xor ((not pi_in(4)(4)(21)) and pi_in(0)(0)(21));
 chi_out(0)(3)(22) <= pi_in(3)(3)(22) xor ((not pi_in(4)(4)(22)) and pi_in(0)(0)(22));
 chi_out(0)(3)(23) <= pi_in(3)(3)(23) xor ((not pi_in(4)(4)(23)) and pi_in(0)(0)(23));
 chi_out(0)(3)(24) <= pi_in(3)(3)(24) xor ((not pi_in(4)(4)(24)) and pi_in(0)(0)(24));
 chi_out(0)(3)(25) <= pi_in(3)(3)(25) xor ((not pi_in(4)(4)(25)) and pi_in(0)(0)(25));
 chi_out(0)(3)(26) <= pi_in(3)(3)(26) xor ((not pi_in(4)(4)(26)) and pi_in(0)(0)(26));
 chi_out(0)(3)(27) <= pi_in(3)(3)(27) xor ((not pi_in(4)(4)(27)) and pi_in(0)(0)(27));
 chi_out(0)(3)(28) <= pi_in(3)(3)(28) xor ((not pi_in(4)(4)(28)) and pi_in(0)(0)(28));
 chi_out(0)(3)(29) <= pi_in(3)(3)(29) xor ((not pi_in(4)(4)(29)) and pi_in(0)(0)(29));
 chi_out(0)(3)(30) <= pi_in(3)(3)(30) xor ((not pi_in(4)(4)(30)) and pi_in(0)(0)(30));
 chi_out(0)(3)(31) <= pi_in(3)(3)(31) xor ((not pi_in(4)(4)(31)) and pi_in(0)(0)(31));
 chi_out(0)(3)(32) <= pi_in(3)(3)(32) xor ((not pi_in(4)(4)(32)) and pi_in(0)(0)(32));
 chi_out(0)(3)(33) <= pi_in(3)(3)(33) xor ((not pi_in(4)(4)(33)) and pi_in(0)(0)(33));
 chi_out(0)(3)(34) <= pi_in(3)(3)(34) xor ((not pi_in(4)(4)(34)) and pi_in(0)(0)(34));
 chi_out(0)(3)(35) <= pi_in(3)(3)(35) xor ((not pi_in(4)(4)(35)) and pi_in(0)(0)(35));
 chi_out(0)(3)(36) <= pi_in(3)(3)(36) xor ((not pi_in(4)(4)(36)) and pi_in(0)(0)(36));
 chi_out(0)(3)(37) <= pi_in(3)(3)(37) xor ((not pi_in(4)(4)(37)) and pi_in(0)(0)(37));
 chi_out(0)(3)(38) <= pi_in(3)(3)(38) xor ((not pi_in(4)(4)(38)) and pi_in(0)(0)(38));
 chi_out(0)(3)(39) <= pi_in(3)(3)(39) xor ((not pi_in(4)(4)(39)) and pi_in(0)(0)(39));
 chi_out(0)(3)(40) <= pi_in(3)(3)(40) xor ((not pi_in(4)(4)(40)) and pi_in(0)(0)(40));
 chi_out(0)(3)(41) <= pi_in(3)(3)(41) xor ((not pi_in(4)(4)(41)) and pi_in(0)(0)(41));
 chi_out(0)(3)(42) <= pi_in(3)(3)(42) xor ((not pi_in(4)(4)(42)) and pi_in(0)(0)(42));
 chi_out(0)(3)(43) <= pi_in(3)(3)(43) xor ((not pi_in(4)(4)(43)) and pi_in(0)(0)(43));
 chi_out(0)(3)(44) <= pi_in(3)(3)(44) xor ((not pi_in(4)(4)(44)) and pi_in(0)(0)(44));
 chi_out(0)(3)(45) <= pi_in(3)(3)(45) xor ((not pi_in(4)(4)(45)) and pi_in(0)(0)(45));
 chi_out(0)(3)(46) <= pi_in(3)(3)(46) xor ((not pi_in(4)(4)(46)) and pi_in(0)(0)(46));
 chi_out(0)(3)(47) <= pi_in(3)(3)(47) xor ((not pi_in(4)(4)(47)) and pi_in(0)(0)(47));
 chi_out(0)(3)(48) <= pi_in(3)(3)(48) xor ((not pi_in(4)(4)(48)) and pi_in(0)(0)(48));
 chi_out(0)(3)(49) <= pi_in(3)(3)(49) xor ((not pi_in(4)(4)(49)) and pi_in(0)(0)(49));
 chi_out(0)(3)(50) <= pi_in(3)(3)(50) xor ((not pi_in(4)(4)(50)) and pi_in(0)(0)(50));
 chi_out(0)(3)(51) <= pi_in(3)(3)(51) xor ((not pi_in(4)(4)(51)) and pi_in(0)(0)(51));
 chi_out(0)(3)(52) <= pi_in(3)(3)(52) xor ((not pi_in(4)(4)(52)) and pi_in(0)(0)(52));
 chi_out(0)(3)(53) <= pi_in(3)(3)(53) xor ((not pi_in(4)(4)(53)) and pi_in(0)(0)(53));
 chi_out(0)(3)(54) <= pi_in(3)(3)(54) xor ((not pi_in(4)(4)(54)) and pi_in(0)(0)(54));
 chi_out(0)(3)(55) <= pi_in(3)(3)(55) xor ((not pi_in(4)(4)(55)) and pi_in(0)(0)(55));
 chi_out(0)(3)(56) <= pi_in(3)(3)(56) xor ((not pi_in(4)(4)(56)) and pi_in(0)(0)(56));
 chi_out(0)(3)(57) <= pi_in(3)(3)(57) xor ((not pi_in(4)(4)(57)) and pi_in(0)(0)(57));
 chi_out(0)(3)(58) <= pi_in(3)(3)(58) xor ((not pi_in(4)(4)(58)) and pi_in(0)(0)(58));
 chi_out(0)(3)(59) <= pi_in(3)(3)(59) xor ((not pi_in(4)(4)(59)) and pi_in(0)(0)(59));
 chi_out(0)(3)(60) <= pi_in(3)(3)(60) xor ((not pi_in(4)(4)(60)) and pi_in(0)(0)(60));
 chi_out(0)(3)(61) <= pi_in(3)(3)(61) xor ((not pi_in(4)(4)(61)) and pi_in(0)(0)(61));
 chi_out(0)(3)(62) <= pi_in(3)(3)(62) xor ((not pi_in(4)(4)(62)) and pi_in(0)(0)(62));
 chi_out(0)(3)(63) <= pi_in(3)(3)(63) xor ((not pi_in(4)(4)(63)) and pi_in(0)(0)(63));
 chi_out(1)(3)(0) <= pi_in(3)(1)(0) xor ((not pi_in(4)(2)(0)) and pi_in(0)(3)(0));
 chi_out(1)(3)(1) <= pi_in(3)(1)(1) xor ((not pi_in(4)(2)(1)) and pi_in(0)(3)(1));
 chi_out(1)(3)(2) <= pi_in(3)(1)(2) xor ((not pi_in(4)(2)(2)) and pi_in(0)(3)(2));
 chi_out(1)(3)(3) <= pi_in(3)(1)(3) xor ((not pi_in(4)(2)(3)) and pi_in(0)(3)(3));
 chi_out(1)(3)(4) <= pi_in(3)(1)(4) xor ((not pi_in(4)(2)(4)) and pi_in(0)(3)(4));
 chi_out(1)(3)(5) <= pi_in(3)(1)(5) xor ((not pi_in(4)(2)(5)) and pi_in(0)(3)(5));
 chi_out(1)(3)(6) <= pi_in(3)(1)(6) xor ((not pi_in(4)(2)(6)) and pi_in(0)(3)(6));
 chi_out(1)(3)(7) <= pi_in(3)(1)(7) xor ((not pi_in(4)(2)(7)) and pi_in(0)(3)(7));
 chi_out(1)(3)(8) <= pi_in(3)(1)(8) xor ((not pi_in(4)(2)(8)) and pi_in(0)(3)(8));
 chi_out(1)(3)(9) <= pi_in(3)(1)(9) xor ((not pi_in(4)(2)(9)) and pi_in(0)(3)(9));
 chi_out(1)(3)(10) <= pi_in(3)(1)(10) xor ((not pi_in(4)(2)(10)) and pi_in(0)(3)(10));
 chi_out(1)(3)(11) <= pi_in(3)(1)(11) xor ((not pi_in(4)(2)(11)) and pi_in(0)(3)(11));
 chi_out(1)(3)(12) <= pi_in(3)(1)(12) xor ((not pi_in(4)(2)(12)) and pi_in(0)(3)(12));
 chi_out(1)(3)(13) <= pi_in(3)(1)(13) xor ((not pi_in(4)(2)(13)) and pi_in(0)(3)(13));
 chi_out(1)(3)(14) <= pi_in(3)(1)(14) xor ((not pi_in(4)(2)(14)) and pi_in(0)(3)(14));
 chi_out(1)(3)(15) <= pi_in(3)(1)(15) xor ((not pi_in(4)(2)(15)) and pi_in(0)(3)(15));
 chi_out(1)(3)(16) <= pi_in(3)(1)(16) xor ((not pi_in(4)(2)(16)) and pi_in(0)(3)(16));
 chi_out(1)(3)(17) <= pi_in(3)(1)(17) xor ((not pi_in(4)(2)(17)) and pi_in(0)(3)(17));
 chi_out(1)(3)(18) <= pi_in(3)(1)(18) xor ((not pi_in(4)(2)(18)) and pi_in(0)(3)(18));
 chi_out(1)(3)(19) <= pi_in(3)(1)(19) xor ((not pi_in(4)(2)(19)) and pi_in(0)(3)(19));
 chi_out(1)(3)(20) <= pi_in(3)(1)(20) xor ((not pi_in(4)(2)(20)) and pi_in(0)(3)(20));
 chi_out(1)(3)(21) <= pi_in(3)(1)(21) xor ((not pi_in(4)(2)(21)) and pi_in(0)(3)(21));
 chi_out(1)(3)(22) <= pi_in(3)(1)(22) xor ((not pi_in(4)(2)(22)) and pi_in(0)(3)(22));
 chi_out(1)(3)(23) <= pi_in(3)(1)(23) xor ((not pi_in(4)(2)(23)) and pi_in(0)(3)(23));
 chi_out(1)(3)(24) <= pi_in(3)(1)(24) xor ((not pi_in(4)(2)(24)) and pi_in(0)(3)(24));
 chi_out(1)(3)(25) <= pi_in(3)(1)(25) xor ((not pi_in(4)(2)(25)) and pi_in(0)(3)(25));
 chi_out(1)(3)(26) <= pi_in(3)(1)(26) xor ((not pi_in(4)(2)(26)) and pi_in(0)(3)(26));
 chi_out(1)(3)(27) <= pi_in(3)(1)(27) xor ((not pi_in(4)(2)(27)) and pi_in(0)(3)(27));
 chi_out(1)(3)(28) <= pi_in(3)(1)(28) xor ((not pi_in(4)(2)(28)) and pi_in(0)(3)(28));
 chi_out(1)(3)(29) <= pi_in(3)(1)(29) xor ((not pi_in(4)(2)(29)) and pi_in(0)(3)(29));
 chi_out(1)(3)(30) <= pi_in(3)(1)(30) xor ((not pi_in(4)(2)(30)) and pi_in(0)(3)(30));
 chi_out(1)(3)(31) <= pi_in(3)(1)(31) xor ((not pi_in(4)(2)(31)) and pi_in(0)(3)(31));
 chi_out(1)(3)(32) <= pi_in(3)(1)(32) xor ((not pi_in(4)(2)(32)) and pi_in(0)(3)(32));
 chi_out(1)(3)(33) <= pi_in(3)(1)(33) xor ((not pi_in(4)(2)(33)) and pi_in(0)(3)(33));
 chi_out(1)(3)(34) <= pi_in(3)(1)(34) xor ((not pi_in(4)(2)(34)) and pi_in(0)(3)(34));
 chi_out(1)(3)(35) <= pi_in(3)(1)(35) xor ((not pi_in(4)(2)(35)) and pi_in(0)(3)(35));
 chi_out(1)(3)(36) <= pi_in(3)(1)(36) xor ((not pi_in(4)(2)(36)) and pi_in(0)(3)(36));
 chi_out(1)(3)(37) <= pi_in(3)(1)(37) xor ((not pi_in(4)(2)(37)) and pi_in(0)(3)(37));
 chi_out(1)(3)(38) <= pi_in(3)(1)(38) xor ((not pi_in(4)(2)(38)) and pi_in(0)(3)(38));
 chi_out(1)(3)(39) <= pi_in(3)(1)(39) xor ((not pi_in(4)(2)(39)) and pi_in(0)(3)(39));
 chi_out(1)(3)(40) <= pi_in(3)(1)(40) xor ((not pi_in(4)(2)(40)) and pi_in(0)(3)(40));
 chi_out(1)(3)(41) <= pi_in(3)(1)(41) xor ((not pi_in(4)(2)(41)) and pi_in(0)(3)(41));
 chi_out(1)(3)(42) <= pi_in(3)(1)(42) xor ((not pi_in(4)(2)(42)) and pi_in(0)(3)(42));
 chi_out(1)(3)(43) <= pi_in(3)(1)(43) xor ((not pi_in(4)(2)(43)) and pi_in(0)(3)(43));
 chi_out(1)(3)(44) <= pi_in(3)(1)(44) xor ((not pi_in(4)(2)(44)) and pi_in(0)(3)(44));
 chi_out(1)(3)(45) <= pi_in(3)(1)(45) xor ((not pi_in(4)(2)(45)) and pi_in(0)(3)(45));
 chi_out(1)(3)(46) <= pi_in(3)(1)(46) xor ((not pi_in(4)(2)(46)) and pi_in(0)(3)(46));
 chi_out(1)(3)(47) <= pi_in(3)(1)(47) xor ((not pi_in(4)(2)(47)) and pi_in(0)(3)(47));
 chi_out(1)(3)(48) <= pi_in(3)(1)(48) xor ((not pi_in(4)(2)(48)) and pi_in(0)(3)(48));
 chi_out(1)(3)(49) <= pi_in(3)(1)(49) xor ((not pi_in(4)(2)(49)) and pi_in(0)(3)(49));
 chi_out(1)(3)(50) <= pi_in(3)(1)(50) xor ((not pi_in(4)(2)(50)) and pi_in(0)(3)(50));
 chi_out(1)(3)(51) <= pi_in(3)(1)(51) xor ((not pi_in(4)(2)(51)) and pi_in(0)(3)(51));
 chi_out(1)(3)(52) <= pi_in(3)(1)(52) xor ((not pi_in(4)(2)(52)) and pi_in(0)(3)(52));
 chi_out(1)(3)(53) <= pi_in(3)(1)(53) xor ((not pi_in(4)(2)(53)) and pi_in(0)(3)(53));
 chi_out(1)(3)(54) <= pi_in(3)(1)(54) xor ((not pi_in(4)(2)(54)) and pi_in(0)(3)(54));
 chi_out(1)(3)(55) <= pi_in(3)(1)(55) xor ((not pi_in(4)(2)(55)) and pi_in(0)(3)(55));
 chi_out(1)(3)(56) <= pi_in(3)(1)(56) xor ((not pi_in(4)(2)(56)) and pi_in(0)(3)(56));
 chi_out(1)(3)(57) <= pi_in(3)(1)(57) xor ((not pi_in(4)(2)(57)) and pi_in(0)(3)(57));
 chi_out(1)(3)(58) <= pi_in(3)(1)(58) xor ((not pi_in(4)(2)(58)) and pi_in(0)(3)(58));
 chi_out(1)(3)(59) <= pi_in(3)(1)(59) xor ((not pi_in(4)(2)(59)) and pi_in(0)(3)(59));
 chi_out(1)(3)(60) <= pi_in(3)(1)(60) xor ((not pi_in(4)(2)(60)) and pi_in(0)(3)(60));
 chi_out(1)(3)(61) <= pi_in(3)(1)(61) xor ((not pi_in(4)(2)(61)) and pi_in(0)(3)(61));
 chi_out(1)(3)(62) <= pi_in(3)(1)(62) xor ((not pi_in(4)(2)(62)) and pi_in(0)(3)(62));
 chi_out(1)(3)(63) <= pi_in(3)(1)(63) xor ((not pi_in(4)(2)(63)) and pi_in(0)(3)(63));
 chi_out(2)(3)(0) <= pi_in(3)(4)(0) xor ((not pi_in(4)(0)(0)) and pi_in(0)(1)(0));
 chi_out(2)(3)(1) <= pi_in(3)(4)(1) xor ((not pi_in(4)(0)(1)) and pi_in(0)(1)(1));
 chi_out(2)(3)(2) <= pi_in(3)(4)(2) xor ((not pi_in(4)(0)(2)) and pi_in(0)(1)(2));
 chi_out(2)(3)(3) <= pi_in(3)(4)(3) xor ((not pi_in(4)(0)(3)) and pi_in(0)(1)(3));
 chi_out(2)(3)(4) <= pi_in(3)(4)(4) xor ((not pi_in(4)(0)(4)) and pi_in(0)(1)(4));
 chi_out(2)(3)(5) <= pi_in(3)(4)(5) xor ((not pi_in(4)(0)(5)) and pi_in(0)(1)(5));
 chi_out(2)(3)(6) <= pi_in(3)(4)(6) xor ((not pi_in(4)(0)(6)) and pi_in(0)(1)(6));
 chi_out(2)(3)(7) <= pi_in(3)(4)(7) xor ((not pi_in(4)(0)(7)) and pi_in(0)(1)(7));
 chi_out(2)(3)(8) <= pi_in(3)(4)(8) xor ((not pi_in(4)(0)(8)) and pi_in(0)(1)(8));
 chi_out(2)(3)(9) <= pi_in(3)(4)(9) xor ((not pi_in(4)(0)(9)) and pi_in(0)(1)(9));
 chi_out(2)(3)(10) <= pi_in(3)(4)(10) xor ((not pi_in(4)(0)(10)) and pi_in(0)(1)(10));
 chi_out(2)(3)(11) <= pi_in(3)(4)(11) xor ((not pi_in(4)(0)(11)) and pi_in(0)(1)(11));
 chi_out(2)(3)(12) <= pi_in(3)(4)(12) xor ((not pi_in(4)(0)(12)) and pi_in(0)(1)(12));
 chi_out(2)(3)(13) <= pi_in(3)(4)(13) xor ((not pi_in(4)(0)(13)) and pi_in(0)(1)(13));
 chi_out(2)(3)(14) <= pi_in(3)(4)(14) xor ((not pi_in(4)(0)(14)) and pi_in(0)(1)(14));
 chi_out(2)(3)(15) <= pi_in(3)(4)(15) xor ((not pi_in(4)(0)(15)) and pi_in(0)(1)(15));
 chi_out(2)(3)(16) <= pi_in(3)(4)(16) xor ((not pi_in(4)(0)(16)) and pi_in(0)(1)(16));
 chi_out(2)(3)(17) <= pi_in(3)(4)(17) xor ((not pi_in(4)(0)(17)) and pi_in(0)(1)(17));
 chi_out(2)(3)(18) <= pi_in(3)(4)(18) xor ((not pi_in(4)(0)(18)) and pi_in(0)(1)(18));
 chi_out(2)(3)(19) <= pi_in(3)(4)(19) xor ((not pi_in(4)(0)(19)) and pi_in(0)(1)(19));
 chi_out(2)(3)(20) <= pi_in(3)(4)(20) xor ((not pi_in(4)(0)(20)) and pi_in(0)(1)(20));
 chi_out(2)(3)(21) <= pi_in(3)(4)(21) xor ((not pi_in(4)(0)(21)) and pi_in(0)(1)(21));
 chi_out(2)(3)(22) <= pi_in(3)(4)(22) xor ((not pi_in(4)(0)(22)) and pi_in(0)(1)(22));
 chi_out(2)(3)(23) <= pi_in(3)(4)(23) xor ((not pi_in(4)(0)(23)) and pi_in(0)(1)(23));
 chi_out(2)(3)(24) <= pi_in(3)(4)(24) xor ((not pi_in(4)(0)(24)) and pi_in(0)(1)(24));
 chi_out(2)(3)(25) <= pi_in(3)(4)(25) xor ((not pi_in(4)(0)(25)) and pi_in(0)(1)(25));
 chi_out(2)(3)(26) <= pi_in(3)(4)(26) xor ((not pi_in(4)(0)(26)) and pi_in(0)(1)(26));
 chi_out(2)(3)(27) <= pi_in(3)(4)(27) xor ((not pi_in(4)(0)(27)) and pi_in(0)(1)(27));
 chi_out(2)(3)(28) <= pi_in(3)(4)(28) xor ((not pi_in(4)(0)(28)) and pi_in(0)(1)(28));
 chi_out(2)(3)(29) <= pi_in(3)(4)(29) xor ((not pi_in(4)(0)(29)) and pi_in(0)(1)(29));
 chi_out(2)(3)(30) <= pi_in(3)(4)(30) xor ((not pi_in(4)(0)(30)) and pi_in(0)(1)(30));
 chi_out(2)(3)(31) <= pi_in(3)(4)(31) xor ((not pi_in(4)(0)(31)) and pi_in(0)(1)(31));
 chi_out(2)(3)(32) <= pi_in(3)(4)(32) xor ((not pi_in(4)(0)(32)) and pi_in(0)(1)(32));
 chi_out(2)(3)(33) <= pi_in(3)(4)(33) xor ((not pi_in(4)(0)(33)) and pi_in(0)(1)(33));
 chi_out(2)(3)(34) <= pi_in(3)(4)(34) xor ((not pi_in(4)(0)(34)) and pi_in(0)(1)(34));
 chi_out(2)(3)(35) <= pi_in(3)(4)(35) xor ((not pi_in(4)(0)(35)) and pi_in(0)(1)(35));
 chi_out(2)(3)(36) <= pi_in(3)(4)(36) xor ((not pi_in(4)(0)(36)) and pi_in(0)(1)(36));
 chi_out(2)(3)(37) <= pi_in(3)(4)(37) xor ((not pi_in(4)(0)(37)) and pi_in(0)(1)(37));
 chi_out(2)(3)(38) <= pi_in(3)(4)(38) xor ((not pi_in(4)(0)(38)) and pi_in(0)(1)(38));
 chi_out(2)(3)(39) <= pi_in(3)(4)(39) xor ((not pi_in(4)(0)(39)) and pi_in(0)(1)(39));
 chi_out(2)(3)(40) <= pi_in(3)(4)(40) xor ((not pi_in(4)(0)(40)) and pi_in(0)(1)(40));
 chi_out(2)(3)(41) <= pi_in(3)(4)(41) xor ((not pi_in(4)(0)(41)) and pi_in(0)(1)(41));
 chi_out(2)(3)(42) <= pi_in(3)(4)(42) xor ((not pi_in(4)(0)(42)) and pi_in(0)(1)(42));
 chi_out(2)(3)(43) <= pi_in(3)(4)(43) xor ((not pi_in(4)(0)(43)) and pi_in(0)(1)(43));
 chi_out(2)(3)(44) <= pi_in(3)(4)(44) xor ((not pi_in(4)(0)(44)) and pi_in(0)(1)(44));
 chi_out(2)(3)(45) <= pi_in(3)(4)(45) xor ((not pi_in(4)(0)(45)) and pi_in(0)(1)(45));
 chi_out(2)(3)(46) <= pi_in(3)(4)(46) xor ((not pi_in(4)(0)(46)) and pi_in(0)(1)(46));
 chi_out(2)(3)(47) <= pi_in(3)(4)(47) xor ((not pi_in(4)(0)(47)) and pi_in(0)(1)(47));
 chi_out(2)(3)(48) <= pi_in(3)(4)(48) xor ((not pi_in(4)(0)(48)) and pi_in(0)(1)(48));
 chi_out(2)(3)(49) <= pi_in(3)(4)(49) xor ((not pi_in(4)(0)(49)) and pi_in(0)(1)(49));
 chi_out(2)(3)(50) <= pi_in(3)(4)(50) xor ((not pi_in(4)(0)(50)) and pi_in(0)(1)(50));
 chi_out(2)(3)(51) <= pi_in(3)(4)(51) xor ((not pi_in(4)(0)(51)) and pi_in(0)(1)(51));
 chi_out(2)(3)(52) <= pi_in(3)(4)(52) xor ((not pi_in(4)(0)(52)) and pi_in(0)(1)(52));
 chi_out(2)(3)(53) <= pi_in(3)(4)(53) xor ((not pi_in(4)(0)(53)) and pi_in(0)(1)(53));
 chi_out(2)(3)(54) <= pi_in(3)(4)(54) xor ((not pi_in(4)(0)(54)) and pi_in(0)(1)(54));
 chi_out(2)(3)(55) <= pi_in(3)(4)(55) xor ((not pi_in(4)(0)(55)) and pi_in(0)(1)(55));
 chi_out(2)(3)(56) <= pi_in(3)(4)(56) xor ((not pi_in(4)(0)(56)) and pi_in(0)(1)(56));
 chi_out(2)(3)(57) <= pi_in(3)(4)(57) xor ((not pi_in(4)(0)(57)) and pi_in(0)(1)(57));
 chi_out(2)(3)(58) <= pi_in(3)(4)(58) xor ((not pi_in(4)(0)(58)) and pi_in(0)(1)(58));
 chi_out(2)(3)(59) <= pi_in(3)(4)(59) xor ((not pi_in(4)(0)(59)) and pi_in(0)(1)(59));
 chi_out(2)(3)(60) <= pi_in(3)(4)(60) xor ((not pi_in(4)(0)(60)) and pi_in(0)(1)(60));
 chi_out(2)(3)(61) <= pi_in(3)(4)(61) xor ((not pi_in(4)(0)(61)) and pi_in(0)(1)(61));
 chi_out(2)(3)(62) <= pi_in(3)(4)(62) xor ((not pi_in(4)(0)(62)) and pi_in(0)(1)(62));
 chi_out(2)(3)(63) <= pi_in(3)(4)(63) xor ((not pi_in(4)(0)(63)) and pi_in(0)(1)(63));
 chi_out(3)(3)(0) <= pi_in(3)(2)(0) xor ((not pi_in(4)(3)(0)) and pi_in(0)(4)(0));
 chi_out(3)(3)(1) <= pi_in(3)(2)(1) xor ((not pi_in(4)(3)(1)) and pi_in(0)(4)(1));
 chi_out(3)(3)(2) <= pi_in(3)(2)(2) xor ((not pi_in(4)(3)(2)) and pi_in(0)(4)(2));
 chi_out(3)(3)(3) <= pi_in(3)(2)(3) xor ((not pi_in(4)(3)(3)) and pi_in(0)(4)(3));
 chi_out(3)(3)(4) <= pi_in(3)(2)(4) xor ((not pi_in(4)(3)(4)) and pi_in(0)(4)(4));
 chi_out(3)(3)(5) <= pi_in(3)(2)(5) xor ((not pi_in(4)(3)(5)) and pi_in(0)(4)(5));
 chi_out(3)(3)(6) <= pi_in(3)(2)(6) xor ((not pi_in(4)(3)(6)) and pi_in(0)(4)(6));
 chi_out(3)(3)(7) <= pi_in(3)(2)(7) xor ((not pi_in(4)(3)(7)) and pi_in(0)(4)(7));
 chi_out(3)(3)(8) <= pi_in(3)(2)(8) xor ((not pi_in(4)(3)(8)) and pi_in(0)(4)(8));
 chi_out(3)(3)(9) <= pi_in(3)(2)(9) xor ((not pi_in(4)(3)(9)) and pi_in(0)(4)(9));
 chi_out(3)(3)(10) <= pi_in(3)(2)(10) xor ((not pi_in(4)(3)(10)) and pi_in(0)(4)(10));
 chi_out(3)(3)(11) <= pi_in(3)(2)(11) xor ((not pi_in(4)(3)(11)) and pi_in(0)(4)(11));
 chi_out(3)(3)(12) <= pi_in(3)(2)(12) xor ((not pi_in(4)(3)(12)) and pi_in(0)(4)(12));
 chi_out(3)(3)(13) <= pi_in(3)(2)(13) xor ((not pi_in(4)(3)(13)) and pi_in(0)(4)(13));
 chi_out(3)(3)(14) <= pi_in(3)(2)(14) xor ((not pi_in(4)(3)(14)) and pi_in(0)(4)(14));
 chi_out(3)(3)(15) <= pi_in(3)(2)(15) xor ((not pi_in(4)(3)(15)) and pi_in(0)(4)(15));
 chi_out(3)(3)(16) <= pi_in(3)(2)(16) xor ((not pi_in(4)(3)(16)) and pi_in(0)(4)(16));
 chi_out(3)(3)(17) <= pi_in(3)(2)(17) xor ((not pi_in(4)(3)(17)) and pi_in(0)(4)(17));
 chi_out(3)(3)(18) <= pi_in(3)(2)(18) xor ((not pi_in(4)(3)(18)) and pi_in(0)(4)(18));
 chi_out(3)(3)(19) <= pi_in(3)(2)(19) xor ((not pi_in(4)(3)(19)) and pi_in(0)(4)(19));
 chi_out(3)(3)(20) <= pi_in(3)(2)(20) xor ((not pi_in(4)(3)(20)) and pi_in(0)(4)(20));
 chi_out(3)(3)(21) <= pi_in(3)(2)(21) xor ((not pi_in(4)(3)(21)) and pi_in(0)(4)(21));
 chi_out(3)(3)(22) <= pi_in(3)(2)(22) xor ((not pi_in(4)(3)(22)) and pi_in(0)(4)(22));
 chi_out(3)(3)(23) <= pi_in(3)(2)(23) xor ((not pi_in(4)(3)(23)) and pi_in(0)(4)(23));
 chi_out(3)(3)(24) <= pi_in(3)(2)(24) xor ((not pi_in(4)(3)(24)) and pi_in(0)(4)(24));
 chi_out(3)(3)(25) <= pi_in(3)(2)(25) xor ((not pi_in(4)(3)(25)) and pi_in(0)(4)(25));
 chi_out(3)(3)(26) <= pi_in(3)(2)(26) xor ((not pi_in(4)(3)(26)) and pi_in(0)(4)(26));
 chi_out(3)(3)(27) <= pi_in(3)(2)(27) xor ((not pi_in(4)(3)(27)) and pi_in(0)(4)(27));
 chi_out(3)(3)(28) <= pi_in(3)(2)(28) xor ((not pi_in(4)(3)(28)) and pi_in(0)(4)(28));
 chi_out(3)(3)(29) <= pi_in(3)(2)(29) xor ((not pi_in(4)(3)(29)) and pi_in(0)(4)(29));
 chi_out(3)(3)(30) <= pi_in(3)(2)(30) xor ((not pi_in(4)(3)(30)) and pi_in(0)(4)(30));
 chi_out(3)(3)(31) <= pi_in(3)(2)(31) xor ((not pi_in(4)(3)(31)) and pi_in(0)(4)(31));
 chi_out(3)(3)(32) <= pi_in(3)(2)(32) xor ((not pi_in(4)(3)(32)) and pi_in(0)(4)(32));
 chi_out(3)(3)(33) <= pi_in(3)(2)(33) xor ((not pi_in(4)(3)(33)) and pi_in(0)(4)(33));
 chi_out(3)(3)(34) <= pi_in(3)(2)(34) xor ((not pi_in(4)(3)(34)) and pi_in(0)(4)(34));
 chi_out(3)(3)(35) <= pi_in(3)(2)(35) xor ((not pi_in(4)(3)(35)) and pi_in(0)(4)(35));
 chi_out(3)(3)(36) <= pi_in(3)(2)(36) xor ((not pi_in(4)(3)(36)) and pi_in(0)(4)(36));
 chi_out(3)(3)(37) <= pi_in(3)(2)(37) xor ((not pi_in(4)(3)(37)) and pi_in(0)(4)(37));
 chi_out(3)(3)(38) <= pi_in(3)(2)(38) xor ((not pi_in(4)(3)(38)) and pi_in(0)(4)(38));
 chi_out(3)(3)(39) <= pi_in(3)(2)(39) xor ((not pi_in(4)(3)(39)) and pi_in(0)(4)(39));
 chi_out(3)(3)(40) <= pi_in(3)(2)(40) xor ((not pi_in(4)(3)(40)) and pi_in(0)(4)(40));
 chi_out(3)(3)(41) <= pi_in(3)(2)(41) xor ((not pi_in(4)(3)(41)) and pi_in(0)(4)(41));
 chi_out(3)(3)(42) <= pi_in(3)(2)(42) xor ((not pi_in(4)(3)(42)) and pi_in(0)(4)(42));
 chi_out(3)(3)(43) <= pi_in(3)(2)(43) xor ((not pi_in(4)(3)(43)) and pi_in(0)(4)(43));
 chi_out(3)(3)(44) <= pi_in(3)(2)(44) xor ((not pi_in(4)(3)(44)) and pi_in(0)(4)(44));
 chi_out(3)(3)(45) <= pi_in(3)(2)(45) xor ((not pi_in(4)(3)(45)) and pi_in(0)(4)(45));
 chi_out(3)(3)(46) <= pi_in(3)(2)(46) xor ((not pi_in(4)(3)(46)) and pi_in(0)(4)(46));
 chi_out(3)(3)(47) <= pi_in(3)(2)(47) xor ((not pi_in(4)(3)(47)) and pi_in(0)(4)(47));
 chi_out(3)(3)(48) <= pi_in(3)(2)(48) xor ((not pi_in(4)(3)(48)) and pi_in(0)(4)(48));
 chi_out(3)(3)(49) <= pi_in(3)(2)(49) xor ((not pi_in(4)(3)(49)) and pi_in(0)(4)(49));
 chi_out(3)(3)(50) <= pi_in(3)(2)(50) xor ((not pi_in(4)(3)(50)) and pi_in(0)(4)(50));
 chi_out(3)(3)(51) <= pi_in(3)(2)(51) xor ((not pi_in(4)(3)(51)) and pi_in(0)(4)(51));
 chi_out(3)(3)(52) <= pi_in(3)(2)(52) xor ((not pi_in(4)(3)(52)) and pi_in(0)(4)(52));
 chi_out(3)(3)(53) <= pi_in(3)(2)(53) xor ((not pi_in(4)(3)(53)) and pi_in(0)(4)(53));
 chi_out(3)(3)(54) <= pi_in(3)(2)(54) xor ((not pi_in(4)(3)(54)) and pi_in(0)(4)(54));
 chi_out(3)(3)(55) <= pi_in(3)(2)(55) xor ((not pi_in(4)(3)(55)) and pi_in(0)(4)(55));
 chi_out(3)(3)(56) <= pi_in(3)(2)(56) xor ((not pi_in(4)(3)(56)) and pi_in(0)(4)(56));
 chi_out(3)(3)(57) <= pi_in(3)(2)(57) xor ((not pi_in(4)(3)(57)) and pi_in(0)(4)(57));
 chi_out(3)(3)(58) <= pi_in(3)(2)(58) xor ((not pi_in(4)(3)(58)) and pi_in(0)(4)(58));
 chi_out(3)(3)(59) <= pi_in(3)(2)(59) xor ((not pi_in(4)(3)(59)) and pi_in(0)(4)(59));
 chi_out(3)(3)(60) <= pi_in(3)(2)(60) xor ((not pi_in(4)(3)(60)) and pi_in(0)(4)(60));
 chi_out(3)(3)(61) <= pi_in(3)(2)(61) xor ((not pi_in(4)(3)(61)) and pi_in(0)(4)(61));
 chi_out(3)(3)(62) <= pi_in(3)(2)(62) xor ((not pi_in(4)(3)(62)) and pi_in(0)(4)(62));
 chi_out(3)(3)(63) <= pi_in(3)(2)(63) xor ((not pi_in(4)(3)(63)) and pi_in(0)(4)(63));
 chi_out(4)(3)(0) <= pi_in(3)(0)(0) xor ((not pi_in(4)(1)(0)) and pi_in(0)(2)(0));
 chi_out(4)(3)(1) <= pi_in(3)(0)(1) xor ((not pi_in(4)(1)(1)) and pi_in(0)(2)(1));
 chi_out(4)(3)(2) <= pi_in(3)(0)(2) xor ((not pi_in(4)(1)(2)) and pi_in(0)(2)(2));
 chi_out(4)(3)(3) <= pi_in(3)(0)(3) xor ((not pi_in(4)(1)(3)) and pi_in(0)(2)(3));
 chi_out(4)(3)(4) <= pi_in(3)(0)(4) xor ((not pi_in(4)(1)(4)) and pi_in(0)(2)(4));
 chi_out(4)(3)(5) <= pi_in(3)(0)(5) xor ((not pi_in(4)(1)(5)) and pi_in(0)(2)(5));
 chi_out(4)(3)(6) <= pi_in(3)(0)(6) xor ((not pi_in(4)(1)(6)) and pi_in(0)(2)(6));
 chi_out(4)(3)(7) <= pi_in(3)(0)(7) xor ((not pi_in(4)(1)(7)) and pi_in(0)(2)(7));
 chi_out(4)(3)(8) <= pi_in(3)(0)(8) xor ((not pi_in(4)(1)(8)) and pi_in(0)(2)(8));
 chi_out(4)(3)(9) <= pi_in(3)(0)(9) xor ((not pi_in(4)(1)(9)) and pi_in(0)(2)(9));
 chi_out(4)(3)(10) <= pi_in(3)(0)(10) xor ((not pi_in(4)(1)(10)) and pi_in(0)(2)(10));
 chi_out(4)(3)(11) <= pi_in(3)(0)(11) xor ((not pi_in(4)(1)(11)) and pi_in(0)(2)(11));
 chi_out(4)(3)(12) <= pi_in(3)(0)(12) xor ((not pi_in(4)(1)(12)) and pi_in(0)(2)(12));
 chi_out(4)(3)(13) <= pi_in(3)(0)(13) xor ((not pi_in(4)(1)(13)) and pi_in(0)(2)(13));
 chi_out(4)(3)(14) <= pi_in(3)(0)(14) xor ((not pi_in(4)(1)(14)) and pi_in(0)(2)(14));
 chi_out(4)(3)(15) <= pi_in(3)(0)(15) xor ((not pi_in(4)(1)(15)) and pi_in(0)(2)(15));
 chi_out(4)(3)(16) <= pi_in(3)(0)(16) xor ((not pi_in(4)(1)(16)) and pi_in(0)(2)(16));
 chi_out(4)(3)(17) <= pi_in(3)(0)(17) xor ((not pi_in(4)(1)(17)) and pi_in(0)(2)(17));
 chi_out(4)(3)(18) <= pi_in(3)(0)(18) xor ((not pi_in(4)(1)(18)) and pi_in(0)(2)(18));
 chi_out(4)(3)(19) <= pi_in(3)(0)(19) xor ((not pi_in(4)(1)(19)) and pi_in(0)(2)(19));
 chi_out(4)(3)(20) <= pi_in(3)(0)(20) xor ((not pi_in(4)(1)(20)) and pi_in(0)(2)(20));
 chi_out(4)(3)(21) <= pi_in(3)(0)(21) xor ((not pi_in(4)(1)(21)) and pi_in(0)(2)(21));
 chi_out(4)(3)(22) <= pi_in(3)(0)(22) xor ((not pi_in(4)(1)(22)) and pi_in(0)(2)(22));
 chi_out(4)(3)(23) <= pi_in(3)(0)(23) xor ((not pi_in(4)(1)(23)) and pi_in(0)(2)(23));
 chi_out(4)(3)(24) <= pi_in(3)(0)(24) xor ((not pi_in(4)(1)(24)) and pi_in(0)(2)(24));
 chi_out(4)(3)(25) <= pi_in(3)(0)(25) xor ((not pi_in(4)(1)(25)) and pi_in(0)(2)(25));
 chi_out(4)(3)(26) <= pi_in(3)(0)(26) xor ((not pi_in(4)(1)(26)) and pi_in(0)(2)(26));
 chi_out(4)(3)(27) <= pi_in(3)(0)(27) xor ((not pi_in(4)(1)(27)) and pi_in(0)(2)(27));
 chi_out(4)(3)(28) <= pi_in(3)(0)(28) xor ((not pi_in(4)(1)(28)) and pi_in(0)(2)(28));
 chi_out(4)(3)(29) <= pi_in(3)(0)(29) xor ((not pi_in(4)(1)(29)) and pi_in(0)(2)(29));
 chi_out(4)(3)(30) <= pi_in(3)(0)(30) xor ((not pi_in(4)(1)(30)) and pi_in(0)(2)(30));
 chi_out(4)(3)(31) <= pi_in(3)(0)(31) xor ((not pi_in(4)(1)(31)) and pi_in(0)(2)(31));
 chi_out(4)(3)(32) <= pi_in(3)(0)(32) xor ((not pi_in(4)(1)(32)) and pi_in(0)(2)(32));
 chi_out(4)(3)(33) <= pi_in(3)(0)(33) xor ((not pi_in(4)(1)(33)) and pi_in(0)(2)(33));
 chi_out(4)(3)(34) <= pi_in(3)(0)(34) xor ((not pi_in(4)(1)(34)) and pi_in(0)(2)(34));
 chi_out(4)(3)(35) <= pi_in(3)(0)(35) xor ((not pi_in(4)(1)(35)) and pi_in(0)(2)(35));
 chi_out(4)(3)(36) <= pi_in(3)(0)(36) xor ((not pi_in(4)(1)(36)) and pi_in(0)(2)(36));
 chi_out(4)(3)(37) <= pi_in(3)(0)(37) xor ((not pi_in(4)(1)(37)) and pi_in(0)(2)(37));
 chi_out(4)(3)(38) <= pi_in(3)(0)(38) xor ((not pi_in(4)(1)(38)) and pi_in(0)(2)(38));
 chi_out(4)(3)(39) <= pi_in(3)(0)(39) xor ((not pi_in(4)(1)(39)) and pi_in(0)(2)(39));
 chi_out(4)(3)(40) <= pi_in(3)(0)(40) xor ((not pi_in(4)(1)(40)) and pi_in(0)(2)(40));
 chi_out(4)(3)(41) <= pi_in(3)(0)(41) xor ((not pi_in(4)(1)(41)) and pi_in(0)(2)(41));
 chi_out(4)(3)(42) <= pi_in(3)(0)(42) xor ((not pi_in(4)(1)(42)) and pi_in(0)(2)(42));
 chi_out(4)(3)(43) <= pi_in(3)(0)(43) xor ((not pi_in(4)(1)(43)) and pi_in(0)(2)(43));
 chi_out(4)(3)(44) <= pi_in(3)(0)(44) xor ((not pi_in(4)(1)(44)) and pi_in(0)(2)(44));
 chi_out(4)(3)(45) <= pi_in(3)(0)(45) xor ((not pi_in(4)(1)(45)) and pi_in(0)(2)(45));
 chi_out(4)(3)(46) <= pi_in(3)(0)(46) xor ((not pi_in(4)(1)(46)) and pi_in(0)(2)(46));
 chi_out(4)(3)(47) <= pi_in(3)(0)(47) xor ((not pi_in(4)(1)(47)) and pi_in(0)(2)(47));
 chi_out(4)(3)(48) <= pi_in(3)(0)(48) xor ((not pi_in(4)(1)(48)) and pi_in(0)(2)(48));
 chi_out(4)(3)(49) <= pi_in(3)(0)(49) xor ((not pi_in(4)(1)(49)) and pi_in(0)(2)(49));
 chi_out(4)(3)(50) <= pi_in(3)(0)(50) xor ((not pi_in(4)(1)(50)) and pi_in(0)(2)(50));
 chi_out(4)(3)(51) <= pi_in(3)(0)(51) xor ((not pi_in(4)(1)(51)) and pi_in(0)(2)(51));
 chi_out(4)(3)(52) <= pi_in(3)(0)(52) xor ((not pi_in(4)(1)(52)) and pi_in(0)(2)(52));
 chi_out(4)(3)(53) <= pi_in(3)(0)(53) xor ((not pi_in(4)(1)(53)) and pi_in(0)(2)(53));
 chi_out(4)(3)(54) <= pi_in(3)(0)(54) xor ((not pi_in(4)(1)(54)) and pi_in(0)(2)(54));
 chi_out(4)(3)(55) <= pi_in(3)(0)(55) xor ((not pi_in(4)(1)(55)) and pi_in(0)(2)(55));
 chi_out(4)(3)(56) <= pi_in(3)(0)(56) xor ((not pi_in(4)(1)(56)) and pi_in(0)(2)(56));
 chi_out(4)(3)(57) <= pi_in(3)(0)(57) xor ((not pi_in(4)(1)(57)) and pi_in(0)(2)(57));
 chi_out(4)(3)(58) <= pi_in(3)(0)(58) xor ((not pi_in(4)(1)(58)) and pi_in(0)(2)(58));
 chi_out(4)(3)(59) <= pi_in(3)(0)(59) xor ((not pi_in(4)(1)(59)) and pi_in(0)(2)(59));
 chi_out(4)(3)(60) <= pi_in(3)(0)(60) xor ((not pi_in(4)(1)(60)) and pi_in(0)(2)(60));
 chi_out(4)(3)(61) <= pi_in(3)(0)(61) xor ((not pi_in(4)(1)(61)) and pi_in(0)(2)(61));
 chi_out(4)(3)(62) <= pi_in(3)(0)(62) xor ((not pi_in(4)(1)(62)) and pi_in(0)(2)(62));
 chi_out(4)(3)(63) <= pi_in(3)(0)(63) xor ((not pi_in(4)(1)(63)) and pi_in(0)(2)(63));
 chi_out(0)(4)(0) <= pi_in(4)(4)(0) xor ((not pi_in(0)(0)(0)) and pi_in(1)(1)(0));
 chi_out(0)(4)(1) <= pi_in(4)(4)(1) xor ((not pi_in(0)(0)(1)) and pi_in(1)(1)(1));
 chi_out(0)(4)(2) <= pi_in(4)(4)(2) xor ((not pi_in(0)(0)(2)) and pi_in(1)(1)(2));
 chi_out(0)(4)(3) <= pi_in(4)(4)(3) xor ((not pi_in(0)(0)(3)) and pi_in(1)(1)(3));
 chi_out(0)(4)(4) <= pi_in(4)(4)(4) xor ((not pi_in(0)(0)(4)) and pi_in(1)(1)(4));
 chi_out(0)(4)(5) <= pi_in(4)(4)(5) xor ((not pi_in(0)(0)(5)) and pi_in(1)(1)(5));
 chi_out(0)(4)(6) <= pi_in(4)(4)(6) xor ((not pi_in(0)(0)(6)) and pi_in(1)(1)(6));
 chi_out(0)(4)(7) <= pi_in(4)(4)(7) xor ((not pi_in(0)(0)(7)) and pi_in(1)(1)(7));
 chi_out(0)(4)(8) <= pi_in(4)(4)(8) xor ((not pi_in(0)(0)(8)) and pi_in(1)(1)(8));
 chi_out(0)(4)(9) <= pi_in(4)(4)(9) xor ((not pi_in(0)(0)(9)) and pi_in(1)(1)(9));
 chi_out(0)(4)(10) <= pi_in(4)(4)(10) xor ((not pi_in(0)(0)(10)) and pi_in(1)(1)(10));
 chi_out(0)(4)(11) <= pi_in(4)(4)(11) xor ((not pi_in(0)(0)(11)) and pi_in(1)(1)(11));
 chi_out(0)(4)(12) <= pi_in(4)(4)(12) xor ((not pi_in(0)(0)(12)) and pi_in(1)(1)(12));
 chi_out(0)(4)(13) <= pi_in(4)(4)(13) xor ((not pi_in(0)(0)(13)) and pi_in(1)(1)(13));
 chi_out(0)(4)(14) <= pi_in(4)(4)(14) xor ((not pi_in(0)(0)(14)) and pi_in(1)(1)(14));
 chi_out(0)(4)(15) <= pi_in(4)(4)(15) xor ((not pi_in(0)(0)(15)) and pi_in(1)(1)(15));
 chi_out(0)(4)(16) <= pi_in(4)(4)(16) xor ((not pi_in(0)(0)(16)) and pi_in(1)(1)(16));
 chi_out(0)(4)(17) <= pi_in(4)(4)(17) xor ((not pi_in(0)(0)(17)) and pi_in(1)(1)(17));
 chi_out(0)(4)(18) <= pi_in(4)(4)(18) xor ((not pi_in(0)(0)(18)) and pi_in(1)(1)(18));
 chi_out(0)(4)(19) <= pi_in(4)(4)(19) xor ((not pi_in(0)(0)(19)) and pi_in(1)(1)(19));
 chi_out(0)(4)(20) <= pi_in(4)(4)(20) xor ((not pi_in(0)(0)(20)) and pi_in(1)(1)(20));
 chi_out(0)(4)(21) <= pi_in(4)(4)(21) xor ((not pi_in(0)(0)(21)) and pi_in(1)(1)(21));
 chi_out(0)(4)(22) <= pi_in(4)(4)(22) xor ((not pi_in(0)(0)(22)) and pi_in(1)(1)(22));
 chi_out(0)(4)(23) <= pi_in(4)(4)(23) xor ((not pi_in(0)(0)(23)) and pi_in(1)(1)(23));
 chi_out(0)(4)(24) <= pi_in(4)(4)(24) xor ((not pi_in(0)(0)(24)) and pi_in(1)(1)(24));
 chi_out(0)(4)(25) <= pi_in(4)(4)(25) xor ((not pi_in(0)(0)(25)) and pi_in(1)(1)(25));
 chi_out(0)(4)(26) <= pi_in(4)(4)(26) xor ((not pi_in(0)(0)(26)) and pi_in(1)(1)(26));
 chi_out(0)(4)(27) <= pi_in(4)(4)(27) xor ((not pi_in(0)(0)(27)) and pi_in(1)(1)(27));
 chi_out(0)(4)(28) <= pi_in(4)(4)(28) xor ((not pi_in(0)(0)(28)) and pi_in(1)(1)(28));
 chi_out(0)(4)(29) <= pi_in(4)(4)(29) xor ((not pi_in(0)(0)(29)) and pi_in(1)(1)(29));
 chi_out(0)(4)(30) <= pi_in(4)(4)(30) xor ((not pi_in(0)(0)(30)) and pi_in(1)(1)(30));
 chi_out(0)(4)(31) <= pi_in(4)(4)(31) xor ((not pi_in(0)(0)(31)) and pi_in(1)(1)(31));
 chi_out(0)(4)(32) <= pi_in(4)(4)(32) xor ((not pi_in(0)(0)(32)) and pi_in(1)(1)(32));
 chi_out(0)(4)(33) <= pi_in(4)(4)(33) xor ((not pi_in(0)(0)(33)) and pi_in(1)(1)(33));
 chi_out(0)(4)(34) <= pi_in(4)(4)(34) xor ((not pi_in(0)(0)(34)) and pi_in(1)(1)(34));
 chi_out(0)(4)(35) <= pi_in(4)(4)(35) xor ((not pi_in(0)(0)(35)) and pi_in(1)(1)(35));
 chi_out(0)(4)(36) <= pi_in(4)(4)(36) xor ((not pi_in(0)(0)(36)) and pi_in(1)(1)(36));
 chi_out(0)(4)(37) <= pi_in(4)(4)(37) xor ((not pi_in(0)(0)(37)) and pi_in(1)(1)(37));
 chi_out(0)(4)(38) <= pi_in(4)(4)(38) xor ((not pi_in(0)(0)(38)) and pi_in(1)(1)(38));
 chi_out(0)(4)(39) <= pi_in(4)(4)(39) xor ((not pi_in(0)(0)(39)) and pi_in(1)(1)(39));
 chi_out(0)(4)(40) <= pi_in(4)(4)(40) xor ((not pi_in(0)(0)(40)) and pi_in(1)(1)(40));
 chi_out(0)(4)(41) <= pi_in(4)(4)(41) xor ((not pi_in(0)(0)(41)) and pi_in(1)(1)(41));
 chi_out(0)(4)(42) <= pi_in(4)(4)(42) xor ((not pi_in(0)(0)(42)) and pi_in(1)(1)(42));
 chi_out(0)(4)(43) <= pi_in(4)(4)(43) xor ((not pi_in(0)(0)(43)) and pi_in(1)(1)(43));
 chi_out(0)(4)(44) <= pi_in(4)(4)(44) xor ((not pi_in(0)(0)(44)) and pi_in(1)(1)(44));
 chi_out(0)(4)(45) <= pi_in(4)(4)(45) xor ((not pi_in(0)(0)(45)) and pi_in(1)(1)(45));
 chi_out(0)(4)(46) <= pi_in(4)(4)(46) xor ((not pi_in(0)(0)(46)) and pi_in(1)(1)(46));
 chi_out(0)(4)(47) <= pi_in(4)(4)(47) xor ((not pi_in(0)(0)(47)) and pi_in(1)(1)(47));
 chi_out(0)(4)(48) <= pi_in(4)(4)(48) xor ((not pi_in(0)(0)(48)) and pi_in(1)(1)(48));
 chi_out(0)(4)(49) <= pi_in(4)(4)(49) xor ((not pi_in(0)(0)(49)) and pi_in(1)(1)(49));
 chi_out(0)(4)(50) <= pi_in(4)(4)(50) xor ((not pi_in(0)(0)(50)) and pi_in(1)(1)(50));
 chi_out(0)(4)(51) <= pi_in(4)(4)(51) xor ((not pi_in(0)(0)(51)) and pi_in(1)(1)(51));
 chi_out(0)(4)(52) <= pi_in(4)(4)(52) xor ((not pi_in(0)(0)(52)) and pi_in(1)(1)(52));
 chi_out(0)(4)(53) <= pi_in(4)(4)(53) xor ((not pi_in(0)(0)(53)) and pi_in(1)(1)(53));
 chi_out(0)(4)(54) <= pi_in(4)(4)(54) xor ((not pi_in(0)(0)(54)) and pi_in(1)(1)(54));
 chi_out(0)(4)(55) <= pi_in(4)(4)(55) xor ((not pi_in(0)(0)(55)) and pi_in(1)(1)(55));
 chi_out(0)(4)(56) <= pi_in(4)(4)(56) xor ((not pi_in(0)(0)(56)) and pi_in(1)(1)(56));
 chi_out(0)(4)(57) <= pi_in(4)(4)(57) xor ((not pi_in(0)(0)(57)) and pi_in(1)(1)(57));
 chi_out(0)(4)(58) <= pi_in(4)(4)(58) xor ((not pi_in(0)(0)(58)) and pi_in(1)(1)(58));
 chi_out(0)(4)(59) <= pi_in(4)(4)(59) xor ((not pi_in(0)(0)(59)) and pi_in(1)(1)(59));
 chi_out(0)(4)(60) <= pi_in(4)(4)(60) xor ((not pi_in(0)(0)(60)) and pi_in(1)(1)(60));
 chi_out(0)(4)(61) <= pi_in(4)(4)(61) xor ((not pi_in(0)(0)(61)) and pi_in(1)(1)(61));
 chi_out(0)(4)(62) <= pi_in(4)(4)(62) xor ((not pi_in(0)(0)(62)) and pi_in(1)(1)(62));
 chi_out(0)(4)(63) <= pi_in(4)(4)(63) xor ((not pi_in(0)(0)(63)) and pi_in(1)(1)(63));
 chi_out(1)(4)(0) <= pi_in(4)(2)(0) xor ((not pi_in(0)(3)(0)) and pi_in(1)(4)(0));
 chi_out(1)(4)(1) <= pi_in(4)(2)(1) xor ((not pi_in(0)(3)(1)) and pi_in(1)(4)(1));
 chi_out(1)(4)(2) <= pi_in(4)(2)(2) xor ((not pi_in(0)(3)(2)) and pi_in(1)(4)(2));
 chi_out(1)(4)(3) <= pi_in(4)(2)(3) xor ((not pi_in(0)(3)(3)) and pi_in(1)(4)(3));
 chi_out(1)(4)(4) <= pi_in(4)(2)(4) xor ((not pi_in(0)(3)(4)) and pi_in(1)(4)(4));
 chi_out(1)(4)(5) <= pi_in(4)(2)(5) xor ((not pi_in(0)(3)(5)) and pi_in(1)(4)(5));
 chi_out(1)(4)(6) <= pi_in(4)(2)(6) xor ((not pi_in(0)(3)(6)) and pi_in(1)(4)(6));
 chi_out(1)(4)(7) <= pi_in(4)(2)(7) xor ((not pi_in(0)(3)(7)) and pi_in(1)(4)(7));
 chi_out(1)(4)(8) <= pi_in(4)(2)(8) xor ((not pi_in(0)(3)(8)) and pi_in(1)(4)(8));
 chi_out(1)(4)(9) <= pi_in(4)(2)(9) xor ((not pi_in(0)(3)(9)) and pi_in(1)(4)(9));
 chi_out(1)(4)(10) <= pi_in(4)(2)(10) xor ((not pi_in(0)(3)(10)) and pi_in(1)(4)(10));
 chi_out(1)(4)(11) <= pi_in(4)(2)(11) xor ((not pi_in(0)(3)(11)) and pi_in(1)(4)(11));
 chi_out(1)(4)(12) <= pi_in(4)(2)(12) xor ((not pi_in(0)(3)(12)) and pi_in(1)(4)(12));
 chi_out(1)(4)(13) <= pi_in(4)(2)(13) xor ((not pi_in(0)(3)(13)) and pi_in(1)(4)(13));
 chi_out(1)(4)(14) <= pi_in(4)(2)(14) xor ((not pi_in(0)(3)(14)) and pi_in(1)(4)(14));
 chi_out(1)(4)(15) <= pi_in(4)(2)(15) xor ((not pi_in(0)(3)(15)) and pi_in(1)(4)(15));
 chi_out(1)(4)(16) <= pi_in(4)(2)(16) xor ((not pi_in(0)(3)(16)) and pi_in(1)(4)(16));
 chi_out(1)(4)(17) <= pi_in(4)(2)(17) xor ((not pi_in(0)(3)(17)) and pi_in(1)(4)(17));
 chi_out(1)(4)(18) <= pi_in(4)(2)(18) xor ((not pi_in(0)(3)(18)) and pi_in(1)(4)(18));
 chi_out(1)(4)(19) <= pi_in(4)(2)(19) xor ((not pi_in(0)(3)(19)) and pi_in(1)(4)(19));
 chi_out(1)(4)(20) <= pi_in(4)(2)(20) xor ((not pi_in(0)(3)(20)) and pi_in(1)(4)(20));
 chi_out(1)(4)(21) <= pi_in(4)(2)(21) xor ((not pi_in(0)(3)(21)) and pi_in(1)(4)(21));
 chi_out(1)(4)(22) <= pi_in(4)(2)(22) xor ((not pi_in(0)(3)(22)) and pi_in(1)(4)(22));
 chi_out(1)(4)(23) <= pi_in(4)(2)(23) xor ((not pi_in(0)(3)(23)) and pi_in(1)(4)(23));
 chi_out(1)(4)(24) <= pi_in(4)(2)(24) xor ((not pi_in(0)(3)(24)) and pi_in(1)(4)(24));
 chi_out(1)(4)(25) <= pi_in(4)(2)(25) xor ((not pi_in(0)(3)(25)) and pi_in(1)(4)(25));
 chi_out(1)(4)(26) <= pi_in(4)(2)(26) xor ((not pi_in(0)(3)(26)) and pi_in(1)(4)(26));
 chi_out(1)(4)(27) <= pi_in(4)(2)(27) xor ((not pi_in(0)(3)(27)) and pi_in(1)(4)(27));
 chi_out(1)(4)(28) <= pi_in(4)(2)(28) xor ((not pi_in(0)(3)(28)) and pi_in(1)(4)(28));
 chi_out(1)(4)(29) <= pi_in(4)(2)(29) xor ((not pi_in(0)(3)(29)) and pi_in(1)(4)(29));
 chi_out(1)(4)(30) <= pi_in(4)(2)(30) xor ((not pi_in(0)(3)(30)) and pi_in(1)(4)(30));
 chi_out(1)(4)(31) <= pi_in(4)(2)(31) xor ((not pi_in(0)(3)(31)) and pi_in(1)(4)(31));
 chi_out(1)(4)(32) <= pi_in(4)(2)(32) xor ((not pi_in(0)(3)(32)) and pi_in(1)(4)(32));
 chi_out(1)(4)(33) <= pi_in(4)(2)(33) xor ((not pi_in(0)(3)(33)) and pi_in(1)(4)(33));
 chi_out(1)(4)(34) <= pi_in(4)(2)(34) xor ((not pi_in(0)(3)(34)) and pi_in(1)(4)(34));
 chi_out(1)(4)(35) <= pi_in(4)(2)(35) xor ((not pi_in(0)(3)(35)) and pi_in(1)(4)(35));
 chi_out(1)(4)(36) <= pi_in(4)(2)(36) xor ((not pi_in(0)(3)(36)) and pi_in(1)(4)(36));
 chi_out(1)(4)(37) <= pi_in(4)(2)(37) xor ((not pi_in(0)(3)(37)) and pi_in(1)(4)(37));
 chi_out(1)(4)(38) <= pi_in(4)(2)(38) xor ((not pi_in(0)(3)(38)) and pi_in(1)(4)(38));
 chi_out(1)(4)(39) <= pi_in(4)(2)(39) xor ((not pi_in(0)(3)(39)) and pi_in(1)(4)(39));
 chi_out(1)(4)(40) <= pi_in(4)(2)(40) xor ((not pi_in(0)(3)(40)) and pi_in(1)(4)(40));
 chi_out(1)(4)(41) <= pi_in(4)(2)(41) xor ((not pi_in(0)(3)(41)) and pi_in(1)(4)(41));
 chi_out(1)(4)(42) <= pi_in(4)(2)(42) xor ((not pi_in(0)(3)(42)) and pi_in(1)(4)(42));
 chi_out(1)(4)(43) <= pi_in(4)(2)(43) xor ((not pi_in(0)(3)(43)) and pi_in(1)(4)(43));
 chi_out(1)(4)(44) <= pi_in(4)(2)(44) xor ((not pi_in(0)(3)(44)) and pi_in(1)(4)(44));
 chi_out(1)(4)(45) <= pi_in(4)(2)(45) xor ((not pi_in(0)(3)(45)) and pi_in(1)(4)(45));
 chi_out(1)(4)(46) <= pi_in(4)(2)(46) xor ((not pi_in(0)(3)(46)) and pi_in(1)(4)(46));
 chi_out(1)(4)(47) <= pi_in(4)(2)(47) xor ((not pi_in(0)(3)(47)) and pi_in(1)(4)(47));
 chi_out(1)(4)(48) <= pi_in(4)(2)(48) xor ((not pi_in(0)(3)(48)) and pi_in(1)(4)(48));
 chi_out(1)(4)(49) <= pi_in(4)(2)(49) xor ((not pi_in(0)(3)(49)) and pi_in(1)(4)(49));
 chi_out(1)(4)(50) <= pi_in(4)(2)(50) xor ((not pi_in(0)(3)(50)) and pi_in(1)(4)(50));
 chi_out(1)(4)(51) <= pi_in(4)(2)(51) xor ((not pi_in(0)(3)(51)) and pi_in(1)(4)(51));
 chi_out(1)(4)(52) <= pi_in(4)(2)(52) xor ((not pi_in(0)(3)(52)) and pi_in(1)(4)(52));
 chi_out(1)(4)(53) <= pi_in(4)(2)(53) xor ((not pi_in(0)(3)(53)) and pi_in(1)(4)(53));
 chi_out(1)(4)(54) <= pi_in(4)(2)(54) xor ((not pi_in(0)(3)(54)) and pi_in(1)(4)(54));
 chi_out(1)(4)(55) <= pi_in(4)(2)(55) xor ((not pi_in(0)(3)(55)) and pi_in(1)(4)(55));
 chi_out(1)(4)(56) <= pi_in(4)(2)(56) xor ((not pi_in(0)(3)(56)) and pi_in(1)(4)(56));
 chi_out(1)(4)(57) <= pi_in(4)(2)(57) xor ((not pi_in(0)(3)(57)) and pi_in(1)(4)(57));
 chi_out(1)(4)(58) <= pi_in(4)(2)(58) xor ((not pi_in(0)(3)(58)) and pi_in(1)(4)(58));
 chi_out(1)(4)(59) <= pi_in(4)(2)(59) xor ((not pi_in(0)(3)(59)) and pi_in(1)(4)(59));
 chi_out(1)(4)(60) <= pi_in(4)(2)(60) xor ((not pi_in(0)(3)(60)) and pi_in(1)(4)(60));
 chi_out(1)(4)(61) <= pi_in(4)(2)(61) xor ((not pi_in(0)(3)(61)) and pi_in(1)(4)(61));
 chi_out(1)(4)(62) <= pi_in(4)(2)(62) xor ((not pi_in(0)(3)(62)) and pi_in(1)(4)(62));
 chi_out(1)(4)(63) <= pi_in(4)(2)(63) xor ((not pi_in(0)(3)(63)) and pi_in(1)(4)(63));
 chi_out(2)(4)(0) <= pi_in(4)(0)(0) xor ((not pi_in(0)(1)(0)) and pi_in(1)(2)(0));
 chi_out(2)(4)(1) <= pi_in(4)(0)(1) xor ((not pi_in(0)(1)(1)) and pi_in(1)(2)(1));
 chi_out(2)(4)(2) <= pi_in(4)(0)(2) xor ((not pi_in(0)(1)(2)) and pi_in(1)(2)(2));
 chi_out(2)(4)(3) <= pi_in(4)(0)(3) xor ((not pi_in(0)(1)(3)) and pi_in(1)(2)(3));
 chi_out(2)(4)(4) <= pi_in(4)(0)(4) xor ((not pi_in(0)(1)(4)) and pi_in(1)(2)(4));
 chi_out(2)(4)(5) <= pi_in(4)(0)(5) xor ((not pi_in(0)(1)(5)) and pi_in(1)(2)(5));
 chi_out(2)(4)(6) <= pi_in(4)(0)(6) xor ((not pi_in(0)(1)(6)) and pi_in(1)(2)(6));
 chi_out(2)(4)(7) <= pi_in(4)(0)(7) xor ((not pi_in(0)(1)(7)) and pi_in(1)(2)(7));
 chi_out(2)(4)(8) <= pi_in(4)(0)(8) xor ((not pi_in(0)(1)(8)) and pi_in(1)(2)(8));
 chi_out(2)(4)(9) <= pi_in(4)(0)(9) xor ((not pi_in(0)(1)(9)) and pi_in(1)(2)(9));
 chi_out(2)(4)(10) <= pi_in(4)(0)(10) xor ((not pi_in(0)(1)(10)) and pi_in(1)(2)(10));
 chi_out(2)(4)(11) <= pi_in(4)(0)(11) xor ((not pi_in(0)(1)(11)) and pi_in(1)(2)(11));
 chi_out(2)(4)(12) <= pi_in(4)(0)(12) xor ((not pi_in(0)(1)(12)) and pi_in(1)(2)(12));
 chi_out(2)(4)(13) <= pi_in(4)(0)(13) xor ((not pi_in(0)(1)(13)) and pi_in(1)(2)(13));
 chi_out(2)(4)(14) <= pi_in(4)(0)(14) xor ((not pi_in(0)(1)(14)) and pi_in(1)(2)(14));
 chi_out(2)(4)(15) <= pi_in(4)(0)(15) xor ((not pi_in(0)(1)(15)) and pi_in(1)(2)(15));
 chi_out(2)(4)(16) <= pi_in(4)(0)(16) xor ((not pi_in(0)(1)(16)) and pi_in(1)(2)(16));
 chi_out(2)(4)(17) <= pi_in(4)(0)(17) xor ((not pi_in(0)(1)(17)) and pi_in(1)(2)(17));
 chi_out(2)(4)(18) <= pi_in(4)(0)(18) xor ((not pi_in(0)(1)(18)) and pi_in(1)(2)(18));
 chi_out(2)(4)(19) <= pi_in(4)(0)(19) xor ((not pi_in(0)(1)(19)) and pi_in(1)(2)(19));
 chi_out(2)(4)(20) <= pi_in(4)(0)(20) xor ((not pi_in(0)(1)(20)) and pi_in(1)(2)(20));
 chi_out(2)(4)(21) <= pi_in(4)(0)(21) xor ((not pi_in(0)(1)(21)) and pi_in(1)(2)(21));
 chi_out(2)(4)(22) <= pi_in(4)(0)(22) xor ((not pi_in(0)(1)(22)) and pi_in(1)(2)(22));
 chi_out(2)(4)(23) <= pi_in(4)(0)(23) xor ((not pi_in(0)(1)(23)) and pi_in(1)(2)(23));
 chi_out(2)(4)(24) <= pi_in(4)(0)(24) xor ((not pi_in(0)(1)(24)) and pi_in(1)(2)(24));
 chi_out(2)(4)(25) <= pi_in(4)(0)(25) xor ((not pi_in(0)(1)(25)) and pi_in(1)(2)(25));
 chi_out(2)(4)(26) <= pi_in(4)(0)(26) xor ((not pi_in(0)(1)(26)) and pi_in(1)(2)(26));
 chi_out(2)(4)(27) <= pi_in(4)(0)(27) xor ((not pi_in(0)(1)(27)) and pi_in(1)(2)(27));
 chi_out(2)(4)(28) <= pi_in(4)(0)(28) xor ((not pi_in(0)(1)(28)) and pi_in(1)(2)(28));
 chi_out(2)(4)(29) <= pi_in(4)(0)(29) xor ((not pi_in(0)(1)(29)) and pi_in(1)(2)(29));
 chi_out(2)(4)(30) <= pi_in(4)(0)(30) xor ((not pi_in(0)(1)(30)) and pi_in(1)(2)(30));
 chi_out(2)(4)(31) <= pi_in(4)(0)(31) xor ((not pi_in(0)(1)(31)) and pi_in(1)(2)(31));
 chi_out(2)(4)(32) <= pi_in(4)(0)(32) xor ((not pi_in(0)(1)(32)) and pi_in(1)(2)(32));
 chi_out(2)(4)(33) <= pi_in(4)(0)(33) xor ((not pi_in(0)(1)(33)) and pi_in(1)(2)(33));
 chi_out(2)(4)(34) <= pi_in(4)(0)(34) xor ((not pi_in(0)(1)(34)) and pi_in(1)(2)(34));
 chi_out(2)(4)(35) <= pi_in(4)(0)(35) xor ((not pi_in(0)(1)(35)) and pi_in(1)(2)(35));
 chi_out(2)(4)(36) <= pi_in(4)(0)(36) xor ((not pi_in(0)(1)(36)) and pi_in(1)(2)(36));
 chi_out(2)(4)(37) <= pi_in(4)(0)(37) xor ((not pi_in(0)(1)(37)) and pi_in(1)(2)(37));
 chi_out(2)(4)(38) <= pi_in(4)(0)(38) xor ((not pi_in(0)(1)(38)) and pi_in(1)(2)(38));
 chi_out(2)(4)(39) <= pi_in(4)(0)(39) xor ((not pi_in(0)(1)(39)) and pi_in(1)(2)(39));
 chi_out(2)(4)(40) <= pi_in(4)(0)(40) xor ((not pi_in(0)(1)(40)) and pi_in(1)(2)(40));
 chi_out(2)(4)(41) <= pi_in(4)(0)(41) xor ((not pi_in(0)(1)(41)) and pi_in(1)(2)(41));
 chi_out(2)(4)(42) <= pi_in(4)(0)(42) xor ((not pi_in(0)(1)(42)) and pi_in(1)(2)(42));
 chi_out(2)(4)(43) <= pi_in(4)(0)(43) xor ((not pi_in(0)(1)(43)) and pi_in(1)(2)(43));
 chi_out(2)(4)(44) <= pi_in(4)(0)(44) xor ((not pi_in(0)(1)(44)) and pi_in(1)(2)(44));
 chi_out(2)(4)(45) <= pi_in(4)(0)(45) xor ((not pi_in(0)(1)(45)) and pi_in(1)(2)(45));
 chi_out(2)(4)(46) <= pi_in(4)(0)(46) xor ((not pi_in(0)(1)(46)) and pi_in(1)(2)(46));
 chi_out(2)(4)(47) <= pi_in(4)(0)(47) xor ((not pi_in(0)(1)(47)) and pi_in(1)(2)(47));
 chi_out(2)(4)(48) <= pi_in(4)(0)(48) xor ((not pi_in(0)(1)(48)) and pi_in(1)(2)(48));
 chi_out(2)(4)(49) <= pi_in(4)(0)(49) xor ((not pi_in(0)(1)(49)) and pi_in(1)(2)(49));
 chi_out(2)(4)(50) <= pi_in(4)(0)(50) xor ((not pi_in(0)(1)(50)) and pi_in(1)(2)(50));
 chi_out(2)(4)(51) <= pi_in(4)(0)(51) xor ((not pi_in(0)(1)(51)) and pi_in(1)(2)(51));
 chi_out(2)(4)(52) <= pi_in(4)(0)(52) xor ((not pi_in(0)(1)(52)) and pi_in(1)(2)(52));
 chi_out(2)(4)(53) <= pi_in(4)(0)(53) xor ((not pi_in(0)(1)(53)) and pi_in(1)(2)(53));
 chi_out(2)(4)(54) <= pi_in(4)(0)(54) xor ((not pi_in(0)(1)(54)) and pi_in(1)(2)(54));
 chi_out(2)(4)(55) <= pi_in(4)(0)(55) xor ((not pi_in(0)(1)(55)) and pi_in(1)(2)(55));
 chi_out(2)(4)(56) <= pi_in(4)(0)(56) xor ((not pi_in(0)(1)(56)) and pi_in(1)(2)(56));
 chi_out(2)(4)(57) <= pi_in(4)(0)(57) xor ((not pi_in(0)(1)(57)) and pi_in(1)(2)(57));
 chi_out(2)(4)(58) <= pi_in(4)(0)(58) xor ((not pi_in(0)(1)(58)) and pi_in(1)(2)(58));
 chi_out(2)(4)(59) <= pi_in(4)(0)(59) xor ((not pi_in(0)(1)(59)) and pi_in(1)(2)(59));
 chi_out(2)(4)(60) <= pi_in(4)(0)(60) xor ((not pi_in(0)(1)(60)) and pi_in(1)(2)(60));
 chi_out(2)(4)(61) <= pi_in(4)(0)(61) xor ((not pi_in(0)(1)(61)) and pi_in(1)(2)(61));
 chi_out(2)(4)(62) <= pi_in(4)(0)(62) xor ((not pi_in(0)(1)(62)) and pi_in(1)(2)(62));
 chi_out(2)(4)(63) <= pi_in(4)(0)(63) xor ((not pi_in(0)(1)(63)) and pi_in(1)(2)(63));
 chi_out(3)(4)(0) <= pi_in(4)(3)(0) xor ((not pi_in(0)(4)(0)) and pi_in(1)(0)(0));
 chi_out(3)(4)(1) <= pi_in(4)(3)(1) xor ((not pi_in(0)(4)(1)) and pi_in(1)(0)(1));
 chi_out(3)(4)(2) <= pi_in(4)(3)(2) xor ((not pi_in(0)(4)(2)) and pi_in(1)(0)(2));
 chi_out(3)(4)(3) <= pi_in(4)(3)(3) xor ((not pi_in(0)(4)(3)) and pi_in(1)(0)(3));
 chi_out(3)(4)(4) <= pi_in(4)(3)(4) xor ((not pi_in(0)(4)(4)) and pi_in(1)(0)(4));
 chi_out(3)(4)(5) <= pi_in(4)(3)(5) xor ((not pi_in(0)(4)(5)) and pi_in(1)(0)(5));
 chi_out(3)(4)(6) <= pi_in(4)(3)(6) xor ((not pi_in(0)(4)(6)) and pi_in(1)(0)(6));
 chi_out(3)(4)(7) <= pi_in(4)(3)(7) xor ((not pi_in(0)(4)(7)) and pi_in(1)(0)(7));
 chi_out(3)(4)(8) <= pi_in(4)(3)(8) xor ((not pi_in(0)(4)(8)) and pi_in(1)(0)(8));
 chi_out(3)(4)(9) <= pi_in(4)(3)(9) xor ((not pi_in(0)(4)(9)) and pi_in(1)(0)(9));
 chi_out(3)(4)(10) <= pi_in(4)(3)(10) xor ((not pi_in(0)(4)(10)) and pi_in(1)(0)(10));
 chi_out(3)(4)(11) <= pi_in(4)(3)(11) xor ((not pi_in(0)(4)(11)) and pi_in(1)(0)(11));
 chi_out(3)(4)(12) <= pi_in(4)(3)(12) xor ((not pi_in(0)(4)(12)) and pi_in(1)(0)(12));
 chi_out(3)(4)(13) <= pi_in(4)(3)(13) xor ((not pi_in(0)(4)(13)) and pi_in(1)(0)(13));
 chi_out(3)(4)(14) <= pi_in(4)(3)(14) xor ((not pi_in(0)(4)(14)) and pi_in(1)(0)(14));
 chi_out(3)(4)(15) <= pi_in(4)(3)(15) xor ((not pi_in(0)(4)(15)) and pi_in(1)(0)(15));
 chi_out(3)(4)(16) <= pi_in(4)(3)(16) xor ((not pi_in(0)(4)(16)) and pi_in(1)(0)(16));
 chi_out(3)(4)(17) <= pi_in(4)(3)(17) xor ((not pi_in(0)(4)(17)) and pi_in(1)(0)(17));
 chi_out(3)(4)(18) <= pi_in(4)(3)(18) xor ((not pi_in(0)(4)(18)) and pi_in(1)(0)(18));
 chi_out(3)(4)(19) <= pi_in(4)(3)(19) xor ((not pi_in(0)(4)(19)) and pi_in(1)(0)(19));
 chi_out(3)(4)(20) <= pi_in(4)(3)(20) xor ((not pi_in(0)(4)(20)) and pi_in(1)(0)(20));
 chi_out(3)(4)(21) <= pi_in(4)(3)(21) xor ((not pi_in(0)(4)(21)) and pi_in(1)(0)(21));
 chi_out(3)(4)(22) <= pi_in(4)(3)(22) xor ((not pi_in(0)(4)(22)) and pi_in(1)(0)(22));
 chi_out(3)(4)(23) <= pi_in(4)(3)(23) xor ((not pi_in(0)(4)(23)) and pi_in(1)(0)(23));
 chi_out(3)(4)(24) <= pi_in(4)(3)(24) xor ((not pi_in(0)(4)(24)) and pi_in(1)(0)(24));
 chi_out(3)(4)(25) <= pi_in(4)(3)(25) xor ((not pi_in(0)(4)(25)) and pi_in(1)(0)(25));
 chi_out(3)(4)(26) <= pi_in(4)(3)(26) xor ((not pi_in(0)(4)(26)) and pi_in(1)(0)(26));
 chi_out(3)(4)(27) <= pi_in(4)(3)(27) xor ((not pi_in(0)(4)(27)) and pi_in(1)(0)(27));
 chi_out(3)(4)(28) <= pi_in(4)(3)(28) xor ((not pi_in(0)(4)(28)) and pi_in(1)(0)(28));
 chi_out(3)(4)(29) <= pi_in(4)(3)(29) xor ((not pi_in(0)(4)(29)) and pi_in(1)(0)(29));
 chi_out(3)(4)(30) <= pi_in(4)(3)(30) xor ((not pi_in(0)(4)(30)) and pi_in(1)(0)(30));
 chi_out(3)(4)(31) <= pi_in(4)(3)(31) xor ((not pi_in(0)(4)(31)) and pi_in(1)(0)(31));
 chi_out(3)(4)(32) <= pi_in(4)(3)(32) xor ((not pi_in(0)(4)(32)) and pi_in(1)(0)(32));
 chi_out(3)(4)(33) <= pi_in(4)(3)(33) xor ((not pi_in(0)(4)(33)) and pi_in(1)(0)(33));
 chi_out(3)(4)(34) <= pi_in(4)(3)(34) xor ((not pi_in(0)(4)(34)) and pi_in(1)(0)(34));
 chi_out(3)(4)(35) <= pi_in(4)(3)(35) xor ((not pi_in(0)(4)(35)) and pi_in(1)(0)(35));
 chi_out(3)(4)(36) <= pi_in(4)(3)(36) xor ((not pi_in(0)(4)(36)) and pi_in(1)(0)(36));
 chi_out(3)(4)(37) <= pi_in(4)(3)(37) xor ((not pi_in(0)(4)(37)) and pi_in(1)(0)(37));
 chi_out(3)(4)(38) <= pi_in(4)(3)(38) xor ((not pi_in(0)(4)(38)) and pi_in(1)(0)(38));
 chi_out(3)(4)(39) <= pi_in(4)(3)(39) xor ((not pi_in(0)(4)(39)) and pi_in(1)(0)(39));
 chi_out(3)(4)(40) <= pi_in(4)(3)(40) xor ((not pi_in(0)(4)(40)) and pi_in(1)(0)(40));
 chi_out(3)(4)(41) <= pi_in(4)(3)(41) xor ((not pi_in(0)(4)(41)) and pi_in(1)(0)(41));
 chi_out(3)(4)(42) <= pi_in(4)(3)(42) xor ((not pi_in(0)(4)(42)) and pi_in(1)(0)(42));
 chi_out(3)(4)(43) <= pi_in(4)(3)(43) xor ((not pi_in(0)(4)(43)) and pi_in(1)(0)(43));
 chi_out(3)(4)(44) <= pi_in(4)(3)(44) xor ((not pi_in(0)(4)(44)) and pi_in(1)(0)(44));
 chi_out(3)(4)(45) <= pi_in(4)(3)(45) xor ((not pi_in(0)(4)(45)) and pi_in(1)(0)(45));
 chi_out(3)(4)(46) <= pi_in(4)(3)(46) xor ((not pi_in(0)(4)(46)) and pi_in(1)(0)(46));
 chi_out(3)(4)(47) <= pi_in(4)(3)(47) xor ((not pi_in(0)(4)(47)) and pi_in(1)(0)(47));
 chi_out(3)(4)(48) <= pi_in(4)(3)(48) xor ((not pi_in(0)(4)(48)) and pi_in(1)(0)(48));
 chi_out(3)(4)(49) <= pi_in(4)(3)(49) xor ((not pi_in(0)(4)(49)) and pi_in(1)(0)(49));
 chi_out(3)(4)(50) <= pi_in(4)(3)(50) xor ((not pi_in(0)(4)(50)) and pi_in(1)(0)(50));
 chi_out(3)(4)(51) <= pi_in(4)(3)(51) xor ((not pi_in(0)(4)(51)) and pi_in(1)(0)(51));
 chi_out(3)(4)(52) <= pi_in(4)(3)(52) xor ((not pi_in(0)(4)(52)) and pi_in(1)(0)(52));
 chi_out(3)(4)(53) <= pi_in(4)(3)(53) xor ((not pi_in(0)(4)(53)) and pi_in(1)(0)(53));
 chi_out(3)(4)(54) <= pi_in(4)(3)(54) xor ((not pi_in(0)(4)(54)) and pi_in(1)(0)(54));
 chi_out(3)(4)(55) <= pi_in(4)(3)(55) xor ((not pi_in(0)(4)(55)) and pi_in(1)(0)(55));
 chi_out(3)(4)(56) <= pi_in(4)(3)(56) xor ((not pi_in(0)(4)(56)) and pi_in(1)(0)(56));
 chi_out(3)(4)(57) <= pi_in(4)(3)(57) xor ((not pi_in(0)(4)(57)) and pi_in(1)(0)(57));
 chi_out(3)(4)(58) <= pi_in(4)(3)(58) xor ((not pi_in(0)(4)(58)) and pi_in(1)(0)(58));
 chi_out(3)(4)(59) <= pi_in(4)(3)(59) xor ((not pi_in(0)(4)(59)) and pi_in(1)(0)(59));
 chi_out(3)(4)(60) <= pi_in(4)(3)(60) xor ((not pi_in(0)(4)(60)) and pi_in(1)(0)(60));
 chi_out(3)(4)(61) <= pi_in(4)(3)(61) xor ((not pi_in(0)(4)(61)) and pi_in(1)(0)(61));
 chi_out(3)(4)(62) <= pi_in(4)(3)(62) xor ((not pi_in(0)(4)(62)) and pi_in(1)(0)(62));
 chi_out(3)(4)(63) <= pi_in(4)(3)(63) xor ((not pi_in(0)(4)(63)) and pi_in(1)(0)(63));
 chi_out(4)(4)(0) <= pi_in(4)(1)(0) xor ((not pi_in(0)(2)(0)) and pi_in(1)(3)(0));
 chi_out(4)(4)(1) <= pi_in(4)(1)(1) xor ((not pi_in(0)(2)(1)) and pi_in(1)(3)(1));
 chi_out(4)(4)(2) <= pi_in(4)(1)(2) xor ((not pi_in(0)(2)(2)) and pi_in(1)(3)(2));
 chi_out(4)(4)(3) <= pi_in(4)(1)(3) xor ((not pi_in(0)(2)(3)) and pi_in(1)(3)(3));
 chi_out(4)(4)(4) <= pi_in(4)(1)(4) xor ((not pi_in(0)(2)(4)) and pi_in(1)(3)(4));
 chi_out(4)(4)(5) <= pi_in(4)(1)(5) xor ((not pi_in(0)(2)(5)) and pi_in(1)(3)(5));
 chi_out(4)(4)(6) <= pi_in(4)(1)(6) xor ((not pi_in(0)(2)(6)) and pi_in(1)(3)(6));
 chi_out(4)(4)(7) <= pi_in(4)(1)(7) xor ((not pi_in(0)(2)(7)) and pi_in(1)(3)(7));
 chi_out(4)(4)(8) <= pi_in(4)(1)(8) xor ((not pi_in(0)(2)(8)) and pi_in(1)(3)(8));
 chi_out(4)(4)(9) <= pi_in(4)(1)(9) xor ((not pi_in(0)(2)(9)) and pi_in(1)(3)(9));
 chi_out(4)(4)(10) <= pi_in(4)(1)(10) xor ((not pi_in(0)(2)(10)) and pi_in(1)(3)(10));
 chi_out(4)(4)(11) <= pi_in(4)(1)(11) xor ((not pi_in(0)(2)(11)) and pi_in(1)(3)(11));
 chi_out(4)(4)(12) <= pi_in(4)(1)(12) xor ((not pi_in(0)(2)(12)) and pi_in(1)(3)(12));
 chi_out(4)(4)(13) <= pi_in(4)(1)(13) xor ((not pi_in(0)(2)(13)) and pi_in(1)(3)(13));
 chi_out(4)(4)(14) <= pi_in(4)(1)(14) xor ((not pi_in(0)(2)(14)) and pi_in(1)(3)(14));
 chi_out(4)(4)(15) <= pi_in(4)(1)(15) xor ((not pi_in(0)(2)(15)) and pi_in(1)(3)(15));
 chi_out(4)(4)(16) <= pi_in(4)(1)(16) xor ((not pi_in(0)(2)(16)) and pi_in(1)(3)(16));
 chi_out(4)(4)(17) <= pi_in(4)(1)(17) xor ((not pi_in(0)(2)(17)) and pi_in(1)(3)(17));
 chi_out(4)(4)(18) <= pi_in(4)(1)(18) xor ((not pi_in(0)(2)(18)) and pi_in(1)(3)(18));
 chi_out(4)(4)(19) <= pi_in(4)(1)(19) xor ((not pi_in(0)(2)(19)) and pi_in(1)(3)(19));
 chi_out(4)(4)(20) <= pi_in(4)(1)(20) xor ((not pi_in(0)(2)(20)) and pi_in(1)(3)(20));
 chi_out(4)(4)(21) <= pi_in(4)(1)(21) xor ((not pi_in(0)(2)(21)) and pi_in(1)(3)(21));
 chi_out(4)(4)(22) <= pi_in(4)(1)(22) xor ((not pi_in(0)(2)(22)) and pi_in(1)(3)(22));
 chi_out(4)(4)(23) <= pi_in(4)(1)(23) xor ((not pi_in(0)(2)(23)) and pi_in(1)(3)(23));
 chi_out(4)(4)(24) <= pi_in(4)(1)(24) xor ((not pi_in(0)(2)(24)) and pi_in(1)(3)(24));
 chi_out(4)(4)(25) <= pi_in(4)(1)(25) xor ((not pi_in(0)(2)(25)) and pi_in(1)(3)(25));
 chi_out(4)(4)(26) <= pi_in(4)(1)(26) xor ((not pi_in(0)(2)(26)) and pi_in(1)(3)(26));
 chi_out(4)(4)(27) <= pi_in(4)(1)(27) xor ((not pi_in(0)(2)(27)) and pi_in(1)(3)(27));
 chi_out(4)(4)(28) <= pi_in(4)(1)(28) xor ((not pi_in(0)(2)(28)) and pi_in(1)(3)(28));
 chi_out(4)(4)(29) <= pi_in(4)(1)(29) xor ((not pi_in(0)(2)(29)) and pi_in(1)(3)(29));
 chi_out(4)(4)(30) <= pi_in(4)(1)(30) xor ((not pi_in(0)(2)(30)) and pi_in(1)(3)(30));
 chi_out(4)(4)(31) <= pi_in(4)(1)(31) xor ((not pi_in(0)(2)(31)) and pi_in(1)(3)(31));
 chi_out(4)(4)(32) <= pi_in(4)(1)(32) xor ((not pi_in(0)(2)(32)) and pi_in(1)(3)(32));
 chi_out(4)(4)(33) <= pi_in(4)(1)(33) xor ((not pi_in(0)(2)(33)) and pi_in(1)(3)(33));
 chi_out(4)(4)(34) <= pi_in(4)(1)(34) xor ((not pi_in(0)(2)(34)) and pi_in(1)(3)(34));
 chi_out(4)(4)(35) <= pi_in(4)(1)(35) xor ((not pi_in(0)(2)(35)) and pi_in(1)(3)(35));
 chi_out(4)(4)(36) <= pi_in(4)(1)(36) xor ((not pi_in(0)(2)(36)) and pi_in(1)(3)(36));
 chi_out(4)(4)(37) <= pi_in(4)(1)(37) xor ((not pi_in(0)(2)(37)) and pi_in(1)(3)(37));
 chi_out(4)(4)(38) <= pi_in(4)(1)(38) xor ((not pi_in(0)(2)(38)) and pi_in(1)(3)(38));
 chi_out(4)(4)(39) <= pi_in(4)(1)(39) xor ((not pi_in(0)(2)(39)) and pi_in(1)(3)(39));
 chi_out(4)(4)(40) <= pi_in(4)(1)(40) xor ((not pi_in(0)(2)(40)) and pi_in(1)(3)(40));
 chi_out(4)(4)(41) <= pi_in(4)(1)(41) xor ((not pi_in(0)(2)(41)) and pi_in(1)(3)(41));
 chi_out(4)(4)(42) <= pi_in(4)(1)(42) xor ((not pi_in(0)(2)(42)) and pi_in(1)(3)(42));
 chi_out(4)(4)(43) <= pi_in(4)(1)(43) xor ((not pi_in(0)(2)(43)) and pi_in(1)(3)(43));
 chi_out(4)(4)(44) <= pi_in(4)(1)(44) xor ((not pi_in(0)(2)(44)) and pi_in(1)(3)(44));
 chi_out(4)(4)(45) <= pi_in(4)(1)(45) xor ((not pi_in(0)(2)(45)) and pi_in(1)(3)(45));
 chi_out(4)(4)(46) <= pi_in(4)(1)(46) xor ((not pi_in(0)(2)(46)) and pi_in(1)(3)(46));
 chi_out(4)(4)(47) <= pi_in(4)(1)(47) xor ((not pi_in(0)(2)(47)) and pi_in(1)(3)(47));
 chi_out(4)(4)(48) <= pi_in(4)(1)(48) xor ((not pi_in(0)(2)(48)) and pi_in(1)(3)(48));
 chi_out(4)(4)(49) <= pi_in(4)(1)(49) xor ((not pi_in(0)(2)(49)) and pi_in(1)(3)(49));
 chi_out(4)(4)(50) <= pi_in(4)(1)(50) xor ((not pi_in(0)(2)(50)) and pi_in(1)(3)(50));
 chi_out(4)(4)(51) <= pi_in(4)(1)(51) xor ((not pi_in(0)(2)(51)) and pi_in(1)(3)(51));
 chi_out(4)(4)(52) <= pi_in(4)(1)(52) xor ((not pi_in(0)(2)(52)) and pi_in(1)(3)(52));
 chi_out(4)(4)(53) <= pi_in(4)(1)(53) xor ((not pi_in(0)(2)(53)) and pi_in(1)(3)(53));
 chi_out(4)(4)(54) <= pi_in(4)(1)(54) xor ((not pi_in(0)(2)(54)) and pi_in(1)(3)(54));
 chi_out(4)(4)(55) <= pi_in(4)(1)(55) xor ((not pi_in(0)(2)(55)) and pi_in(1)(3)(55));
 chi_out(4)(4)(56) <= pi_in(4)(1)(56) xor ((not pi_in(0)(2)(56)) and pi_in(1)(3)(56));
 chi_out(4)(4)(57) <= pi_in(4)(1)(57) xor ((not pi_in(0)(2)(57)) and pi_in(1)(3)(57));
 chi_out(4)(4)(58) <= pi_in(4)(1)(58) xor ((not pi_in(0)(2)(58)) and pi_in(1)(3)(58));
 chi_out(4)(4)(59) <= pi_in(4)(1)(59) xor ((not pi_in(0)(2)(59)) and pi_in(1)(3)(59));
 chi_out(4)(4)(60) <= pi_in(4)(1)(60) xor ((not pi_in(0)(2)(60)) and pi_in(1)(3)(60));
 chi_out(4)(4)(61) <= pi_in(4)(1)(61) xor ((not pi_in(0)(2)(61)) and pi_in(1)(3)(61));
 chi_out(4)(4)(62) <= pi_in(4)(1)(62) xor ((not pi_in(0)(2)(62)) and pi_in(1)(3)(62));
 chi_out(4)(4)(63) <= pi_in(4)(1)(63) xor ((not pi_in(0)(2)(63)) and pi_in(1)(3)(63));
 



    rho_pi_chi_out<= chi_out;

end architecture RTL;
